magic
tech scmos
timestamp 1635828931
<< nwell >>
rect 27 20 57 36
<< polysilicon >>
rect 34 28 36 30
rect 38 28 40 30
rect 34 20 36 22
rect 35 16 36 20
rect 38 20 40 22
rect 38 19 50 20
rect 38 18 49 19
rect 34 14 40 16
rect 38 12 40 14
rect 48 15 49 18
rect 48 12 50 15
rect 38 7 40 9
rect 48 7 50 9
<< ndiffusion >>
rect 37 9 38 12
rect 40 9 42 12
rect 46 9 48 12
rect 50 9 51 12
<< pdiffusion >>
rect 33 25 34 28
rect 30 22 34 25
rect 36 22 38 28
rect 40 26 45 28
rect 40 22 42 26
<< metal1 >>
rect 31 33 35 36
rect 39 33 43 36
rect 47 33 51 36
rect 55 33 57 36
rect 27 32 57 33
rect 29 29 33 32
rect 46 22 48 26
rect 29 16 31 19
rect 42 12 46 22
rect 53 15 55 18
rect 33 4 37 8
rect 51 4 55 8
rect 27 0 32 3
rect 36 3 37 4
rect 36 0 40 3
rect 44 0 48 3
rect 52 3 55 4
rect 52 0 57 3
<< metal2 >>
rect 52 22 53 26
<< ntransistor >>
rect 38 9 40 12
rect 48 9 50 12
<< ptransistor >>
rect 34 22 36 28
rect 38 22 40 28
<< polycontact >>
rect 31 16 35 20
rect 49 15 53 19
<< ndcontact >>
rect 33 8 37 12
rect 42 8 46 12
rect 51 8 55 12
<< pdcontact >>
rect 29 25 33 29
rect 42 22 46 26
<< m2contact >>
rect 48 22 52 26
<< psubstratepcontact >>
rect 32 0 36 4
rect 40 0 44 4
rect 48 0 52 4
<< nsubstratencontact >>
rect 27 33 31 37
rect 35 33 39 37
rect 43 33 47 37
rect 51 33 55 37
<< labels >>
rlabel metal1 41 34 41 34 5 V_DD
rlabel metal1 39 1 39 1 1 gnd
rlabel metal1 54 17 54 17 7 B
rlabel metal1 30 18 30 18 3 A
rlabel m2contact 52 24 52 24 7 out
rlabel pdiffusion 37 25 37 25 1 pun_mid_node
<< end >>
