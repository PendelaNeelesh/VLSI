*pseudo nmos load
.include ./cmos_include.txt

m2 out 0 vdd vdd cmosp l=1u w=4u
m1 out in 0 0 cmosn l=1u w=2u

Vdd vdd 0 5
V_in in 0 pulse(0 5 0.1n 0.1n 0.1n 2n 4n)

.dc V_in 0 5 0.1

.control
    foreach wid in 1u 10u 100u
    alter @m1 w=$wid
    run
    plot out
    end
.endc

.end
