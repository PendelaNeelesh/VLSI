* SPICE3 file created from cmos_nand_layout.ext - technology: scmos

.model pfet pmos level=3 version=3.3.0
.model nfet nmos level=3 version=3.3.0

.option scale=1u

M1000 pdn_a_b A gnd Gnd nfet w=3 l=2
+  ad=12 pd=14 as=22 ps=20
M1001 out A V_DD V_DD pfet w=6 l=2
+  ad=48 pd=28 as=68 ps=48
M1002 V_DD B out V_DD pfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 out B pdn_a_b Gnd nfet w=3 l=2
+  ad=22 pd=20 as=0 ps=0
C0 A V_DD 2.07fF
C1 gnd Gnd 4.18fF
C2 out Gnd 3.20fF
C3 B Gnd 7.04fF
C4 A Gnd 5.45fF

V_A A gnd pulse(0 5 0.1n 0.1n 0.1n 4n 8n)
V_B B gnd pulse(0 5 0.1n 0.1n 0.1n 2n 4n)
v_dd V_DD gnd 5

.control
	tran 0.1n 16n
	setplot tran1
	plot A B out
.endc

.end
