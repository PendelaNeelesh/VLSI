* SPICE3 file created from cmos_nor_layout.ext - technology: scmos

.model pfet pmos level=3 version=3.3.0
.model nfet nmos level=3 version=3.3.0

.option scale=1u

M1000 pun_mid_node A V_DD V_DD pfet w=6 l=2
+  ad=12 pd=16 as=31 ps=24
M1001 gnd B out Gnd nfet w=3 l=2
+  ad=38 pd=36 as=28 ps=24
M1002 out A gnd Gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 out B pun_mid_node V_DD pfet w=6 l=2
+  ad=34 pd=24 as=0 ps=0
C0 V_DD B 2.23fF
C1 gnd Gnd 4.23fF
C2 B Gnd 5.53fF
C3 A Gnd 4.66fF


V_A A gnd pulse(0 5 0.1n 0.1n 0.1n 4n 8n)
V_B B gnd pulse(0 5 0.1n 0.1n 0.1n 2n 4n)
v_dd V_DD gnd 5

.control
	tran 0.1n 16n
	setplot tran1
	plot A B out
.endc

.end
