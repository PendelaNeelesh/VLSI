magic
tech scmos
timestamp 1635954421
<< ab >>
rect -56 23 0 95
rect 6 59 46 95
rect 50 59 82 95
rect 6 55 44 59
rect 6 23 46 55
rect 50 54 52 55
rect 56 54 82 59
rect 50 23 82 54
rect -56 -67 0 5
rect 4 -67 44 5
<< nwell >>
rect -61 55 82 100
rect -61 -72 49 -27
<< pwell >>
rect -61 23 82 55
rect -61 -27 49 5
<< poly >>
rect -31 89 -29 93
rect -21 89 -19 93
rect -11 89 -9 93
rect 15 89 17 93
rect 25 89 27 93
rect 35 89 37 93
rect 61 89 63 93
rect 68 89 70 93
rect -41 81 -39 85
rect 15 66 17 70
rect 11 64 17 66
rect 11 62 13 64
rect 15 62 17 64
rect -41 58 -39 61
rect -31 58 -29 61
rect -21 58 -19 61
rect -11 58 -9 61
rect 11 60 17 62
rect -41 56 -9 58
rect -41 54 -39 56
rect -37 54 -31 56
rect -29 54 -27 56
rect -41 52 -27 54
rect -41 49 -39 52
rect -31 49 -29 52
rect -21 49 -19 56
rect -11 49 -9 56
rect 15 49 17 60
rect 25 58 27 70
rect 35 58 37 61
rect 21 56 27 58
rect 21 54 23 56
rect 25 54 27 56
rect 21 52 27 54
rect 31 56 37 58
rect 31 54 33 56
rect 35 54 37 56
rect 61 55 63 61
rect 68 58 70 61
rect 31 52 37 54
rect 22 49 24 52
rect 35 49 37 52
rect 57 53 63 55
rect 57 51 59 53
rect 61 51 63 53
rect 67 56 73 58
rect 67 54 69 56
rect 71 54 73 56
rect 67 52 73 54
rect 57 49 63 51
rect -11 35 -9 40
rect 15 31 17 36
rect 22 31 24 36
rect 59 46 61 49
rect 70 43 72 52
rect -41 25 -39 29
rect -31 25 -29 29
rect -21 25 -19 29
rect 35 30 37 35
rect 59 34 61 38
rect 70 30 72 35
rect -41 -1 -39 3
rect -31 -1 -29 3
rect -21 -1 -19 3
rect -11 -12 -9 -7
rect 13 -8 15 -3
rect 20 -8 22 -3
rect 33 -7 35 -2
rect -41 -24 -39 -21
rect -31 -24 -29 -21
rect -41 -26 -27 -24
rect -41 -28 -39 -26
rect -37 -28 -31 -26
rect -29 -28 -27 -26
rect -21 -28 -19 -21
rect -11 -28 -9 -21
rect -41 -30 -9 -28
rect -41 -33 -39 -30
rect -31 -33 -29 -30
rect -21 -33 -19 -30
rect -11 -33 -9 -30
rect 13 -32 15 -21
rect 20 -24 22 -21
rect 33 -24 35 -21
rect 19 -26 25 -24
rect 19 -28 21 -26
rect 23 -28 25 -26
rect 19 -30 25 -28
rect 29 -26 35 -24
rect 29 -28 31 -26
rect 33 -28 35 -26
rect 29 -30 35 -28
rect -41 -57 -39 -53
rect 9 -34 15 -32
rect 9 -36 11 -34
rect 13 -36 15 -34
rect 9 -38 15 -36
rect 13 -42 15 -38
rect 23 -42 25 -30
rect 33 -33 35 -30
rect -31 -65 -29 -61
rect -21 -65 -19 -61
rect -11 -65 -9 -61
rect 13 -65 15 -61
rect 23 -65 25 -61
rect 33 -65 35 -61
<< ndif >>
rect -49 40 -41 49
rect -49 38 -47 40
rect -45 38 -41 40
rect -49 33 -41 38
rect -49 31 -47 33
rect -45 31 -41 33
rect -49 29 -41 31
rect -39 47 -31 49
rect -39 45 -36 47
rect -34 45 -31 47
rect -39 40 -31 45
rect -39 38 -36 40
rect -34 38 -31 40
rect -39 29 -31 38
rect -29 40 -21 49
rect -29 38 -26 40
rect -24 38 -21 40
rect -29 33 -21 38
rect -29 31 -26 33
rect -24 31 -21 33
rect -29 29 -21 31
rect -19 47 -11 49
rect -19 45 -16 47
rect -14 45 -11 47
rect -19 40 -11 45
rect -9 44 -2 49
rect -9 42 -6 44
rect -4 42 -2 44
rect 10 42 15 49
rect -9 40 -2 42
rect 8 40 15 42
rect -19 29 -14 40
rect 8 38 10 40
rect 12 38 15 40
rect 8 36 15 38
rect 17 36 22 49
rect 24 36 35 49
rect 26 35 35 36
rect 37 47 44 49
rect 37 45 40 47
rect 42 45 44 47
rect 37 39 44 45
rect 37 37 40 39
rect 42 37 44 39
rect 52 42 59 46
rect 52 40 54 42
rect 56 40 59 42
rect 52 38 59 40
rect 61 43 66 46
rect 61 39 70 43
rect 61 38 65 39
rect 37 35 44 37
rect 26 30 33 35
rect 63 37 65 38
rect 67 37 70 39
rect 63 35 70 37
rect 72 35 80 43
rect 74 30 80 35
rect 26 28 29 30
rect 31 28 33 30
rect 26 26 33 28
rect 74 28 76 30
rect 78 28 80 30
rect 74 26 80 28
rect -49 -3 -41 -1
rect -49 -5 -47 -3
rect -45 -5 -41 -3
rect -49 -10 -41 -5
rect -49 -12 -47 -10
rect -45 -12 -41 -10
rect -49 -21 -41 -12
rect -39 -10 -31 -1
rect -39 -12 -36 -10
rect -34 -12 -31 -10
rect -39 -17 -31 -12
rect -39 -19 -36 -17
rect -34 -19 -31 -17
rect -39 -21 -31 -19
rect -29 -3 -21 -1
rect -29 -5 -26 -3
rect -24 -5 -21 -3
rect -29 -10 -21 -5
rect -29 -12 -26 -10
rect -24 -12 -21 -10
rect -29 -21 -21 -12
rect -19 -12 -14 -1
rect 24 0 31 2
rect 24 -2 27 0
rect 29 -2 31 0
rect 24 -7 31 -2
rect 24 -8 33 -7
rect 6 -10 13 -8
rect 6 -12 8 -10
rect 10 -12 13 -10
rect -19 -17 -11 -12
rect -19 -19 -16 -17
rect -14 -19 -11 -17
rect -19 -21 -11 -19
rect -9 -14 -2 -12
rect 6 -14 13 -12
rect -9 -16 -6 -14
rect -4 -16 -2 -14
rect -9 -21 -2 -16
rect 8 -21 13 -14
rect 15 -21 20 -8
rect 22 -21 33 -8
rect 35 -9 42 -7
rect 35 -11 38 -9
rect 40 -11 42 -9
rect 35 -17 42 -11
rect 35 -19 38 -17
rect 40 -19 42 -17
rect 35 -21 42 -19
<< pdif >>
rect -36 81 -31 89
rect -48 79 -41 81
rect -48 77 -46 79
rect -44 77 -41 79
rect -48 72 -41 77
rect -48 70 -46 72
rect -44 70 -41 72
rect -48 61 -41 70
rect -39 72 -31 81
rect -39 70 -36 72
rect -34 70 -31 72
rect -39 65 -31 70
rect -39 63 -36 65
rect -34 63 -31 65
rect -39 61 -31 63
rect -29 87 -21 89
rect -29 85 -26 87
rect -24 85 -21 87
rect -29 79 -21 85
rect -29 77 -26 79
rect -24 77 -21 79
rect -29 61 -21 77
rect -19 72 -11 89
rect -19 70 -16 72
rect -14 70 -11 72
rect -19 65 -11 70
rect -19 63 -16 65
rect -14 63 -11 65
rect -19 61 -11 63
rect -9 87 -2 89
rect -9 85 -6 87
rect -4 85 -2 87
rect -9 80 -2 85
rect -9 78 -6 80
rect -4 78 -2 80
rect -9 61 -2 78
rect 8 87 15 89
rect 8 85 10 87
rect 12 85 15 87
rect 8 80 15 85
rect 8 78 10 80
rect 12 78 15 80
rect 8 70 15 78
rect 17 81 25 89
rect 17 79 20 81
rect 22 79 25 81
rect 17 74 25 79
rect 17 72 20 74
rect 22 72 25 74
rect 17 70 25 72
rect 27 87 35 89
rect 27 85 30 87
rect 32 85 35 87
rect 27 80 35 85
rect 27 78 30 80
rect 32 78 35 80
rect 27 70 35 78
rect 29 61 35 70
rect 37 82 42 89
rect 52 87 61 89
rect 52 85 54 87
rect 56 85 61 87
rect 37 80 44 82
rect 37 78 40 80
rect 42 78 44 80
rect 37 73 44 78
rect 37 71 40 73
rect 42 71 44 73
rect 37 69 44 71
rect 52 80 61 85
rect 52 78 54 80
rect 56 78 61 80
rect 37 61 42 69
rect 52 61 61 78
rect 63 61 68 89
rect 70 82 75 89
rect 70 80 77 82
rect 70 78 73 80
rect 75 78 77 80
rect 70 73 77 78
rect 70 71 73 73
rect 75 71 77 73
rect 70 69 77 71
rect 70 61 75 69
rect -48 -42 -41 -33
rect -48 -44 -46 -42
rect -44 -44 -41 -42
rect -48 -49 -41 -44
rect -48 -51 -46 -49
rect -44 -51 -41 -49
rect -48 -53 -41 -51
rect -39 -35 -31 -33
rect -39 -37 -36 -35
rect -34 -37 -31 -35
rect -39 -42 -31 -37
rect -39 -44 -36 -42
rect -34 -44 -31 -42
rect -39 -53 -31 -44
rect -36 -61 -31 -53
rect -29 -49 -21 -33
rect -29 -51 -26 -49
rect -24 -51 -21 -49
rect -29 -57 -21 -51
rect -29 -59 -26 -57
rect -24 -59 -21 -57
rect -29 -61 -21 -59
rect -19 -35 -11 -33
rect -19 -37 -16 -35
rect -14 -37 -11 -35
rect -19 -42 -11 -37
rect -19 -44 -16 -42
rect -14 -44 -11 -42
rect -19 -61 -11 -44
rect -9 -50 -2 -33
rect 27 -42 33 -33
rect -9 -52 -6 -50
rect -4 -52 -2 -50
rect -9 -57 -2 -52
rect -9 -59 -6 -57
rect -4 -59 -2 -57
rect -9 -61 -2 -59
rect 6 -50 13 -42
rect 6 -52 8 -50
rect 10 -52 13 -50
rect 6 -57 13 -52
rect 6 -59 8 -57
rect 10 -59 13 -57
rect 6 -61 13 -59
rect 15 -44 23 -42
rect 15 -46 18 -44
rect 20 -46 23 -44
rect 15 -51 23 -46
rect 15 -53 18 -51
rect 20 -53 23 -51
rect 15 -61 23 -53
rect 25 -50 33 -42
rect 25 -52 28 -50
rect 30 -52 33 -50
rect 25 -57 33 -52
rect 25 -59 28 -57
rect 30 -59 33 -57
rect 25 -61 33 -59
rect 35 -41 40 -33
rect 35 -43 42 -41
rect 35 -45 38 -43
rect 40 -45 42 -43
rect 35 -50 42 -45
rect 35 -52 38 -50
rect 40 -52 42 -50
rect 35 -54 42 -52
rect 35 -61 40 -54
<< alu1 >>
rect -74 90 82 95
rect -74 88 -51 90
rect -49 88 82 90
rect -74 87 82 88
rect -74 -59 -66 87
rect 39 80 44 82
rect 39 78 40 80
rect 42 78 44 80
rect -38 72 -33 74
rect -38 70 -36 72
rect -34 70 -33 72
rect -46 58 -42 66
rect -38 65 -33 70
rect -14 65 -10 66
rect 8 65 12 74
rect 39 73 44 78
rect 71 80 77 81
rect 71 78 73 80
rect 75 78 77 80
rect 39 71 40 73
rect 42 71 44 73
rect 39 69 44 71
rect 71 74 77 78
rect 71 73 80 74
rect 71 71 73 73
rect 75 71 80 73
rect 71 70 80 71
rect 40 66 44 69
rect -38 63 -36 65
rect -34 63 -16 65
rect -14 64 21 65
rect -14 63 13 64
rect -38 62 13 63
rect 15 62 21 64
rect -38 61 21 62
rect -61 57 -42 58
rect -61 55 -59 57
rect -57 56 -25 57
rect -57 55 -39 56
rect -61 54 -39 55
rect -37 54 -31 56
rect -29 54 -25 56
rect -61 53 -25 54
rect -14 49 -10 61
rect -39 47 -10 49
rect -39 45 -36 47
rect -34 45 -16 47
rect -14 45 -10 47
rect 15 56 29 57
rect 15 54 23 56
rect 25 54 29 56
rect 15 53 29 54
rect 15 47 20 53
rect 40 62 64 66
rect 40 61 72 62
rect -39 40 -33 45
rect -18 44 -10 45
rect 15 45 17 47
rect 19 45 20 47
rect 15 44 20 45
rect -39 38 -36 40
rect -34 38 -33 40
rect -39 36 -33 38
rect 40 47 44 61
rect 60 58 72 61
rect 68 56 72 58
rect 68 54 69 56
rect 71 54 72 56
rect 48 53 64 54
rect 48 51 49 53
rect 51 51 59 53
rect 61 51 64 53
rect 68 52 72 54
rect 48 50 64 51
rect 42 45 44 47
rect 40 42 44 45
rect 60 44 64 50
rect 32 39 44 42
rect 32 37 40 39
rect 42 37 44 39
rect 32 36 44 37
rect 76 42 80 70
rect 68 40 80 42
rect 63 39 80 40
rect 63 37 65 39
rect 67 37 80 39
rect 63 36 80 37
rect -58 30 82 31
rect -58 28 -7 30
rect -5 28 29 30
rect 31 28 55 30
rect 57 28 76 30
rect 78 28 82 30
rect -58 23 82 28
rect -58 5 -46 23
rect -58 0 46 5
rect -58 -2 -7 0
rect -5 -2 27 0
rect 29 -2 46 0
rect -58 -3 46 -2
rect -39 -10 -33 -8
rect -39 -12 -36 -10
rect -34 -12 -33 -10
rect -39 -17 -33 -12
rect 30 -9 42 -8
rect -18 -17 -10 -16
rect -39 -19 -36 -17
rect -34 -19 -16 -17
rect -14 -19 -10 -17
rect -39 -21 -10 -19
rect -50 -26 -25 -25
rect -50 -28 -49 -26
rect -47 -28 -39 -26
rect -37 -28 -31 -26
rect -29 -28 -25 -26
rect -50 -29 -25 -28
rect -46 -38 -42 -29
rect -14 -33 -10 -21
rect 13 -25 18 -16
rect 30 -11 38 -9
rect 40 -11 42 -9
rect 30 -14 42 -11
rect 38 -17 42 -14
rect 40 -19 42 -17
rect 0 -26 27 -25
rect 0 -28 2 -26
rect 4 -28 21 -26
rect 23 -28 27 -26
rect 0 -29 27 -28
rect -38 -34 19 -33
rect -38 -35 11 -34
rect -38 -37 -36 -35
rect -34 -37 -16 -35
rect -14 -36 11 -35
rect 13 -36 19 -34
rect -14 -37 19 -36
rect 38 -28 42 -19
rect 38 -30 39 -28
rect 41 -30 42 -28
rect -38 -42 -33 -37
rect -38 -44 -36 -42
rect -34 -44 -33 -42
rect -38 -46 -33 -44
rect -14 -38 -10 -37
rect 6 -46 10 -37
rect 38 -41 42 -30
rect 37 -43 42 -41
rect 37 -45 38 -43
rect 40 -45 42 -43
rect 37 -50 42 -45
rect 37 -52 38 -50
rect 40 -52 42 -50
rect 37 -54 42 -52
rect -74 -60 46 -59
rect -74 -62 -51 -60
rect -49 -62 46 -60
rect -74 -67 46 -62
<< alu2 >>
rect -61 57 -55 58
rect -61 55 -59 57
rect -57 55 -55 57
rect -61 23 -55 55
rect 47 53 52 54
rect 47 51 49 53
rect 51 51 52 53
rect 47 50 52 51
rect 15 47 20 48
rect 15 45 17 47
rect 19 45 20 47
rect 15 44 20 45
rect -61 18 6 23
rect -50 -26 -46 -25
rect -50 -28 -49 -26
rect -47 -28 -46 -26
rect -50 -29 -46 -28
rect 0 -26 6 18
rect 0 -28 2 -26
rect 4 -28 6 -26
rect 0 -29 6 -28
rect 38 -28 46 -27
rect 38 -30 39 -28
rect 41 -30 46 -28
rect 38 -31 46 -30
<< alu3 >>
rect 47 53 52 54
rect 47 51 49 53
rect 51 51 52 53
rect 47 50 52 51
rect 15 47 20 48
rect 15 45 17 47
rect 19 45 20 47
rect 15 10 20 45
rect -61 5 20 10
rect -61 -25 -57 5
rect -61 -26 -46 -25
rect -61 -28 -49 -26
rect -47 -28 -46 -26
rect -61 -29 -46 -28
rect 38 -28 46 -27
rect 38 -30 39 -28
rect 41 -30 46 -28
rect 38 -31 46 -30
<< alu4 >>
rect 44 53 52 54
rect 44 51 49 53
rect 51 51 52 53
rect 44 50 52 51
rect 44 43 50 50
rect 43 42 50 43
rect 43 -23 49 42
rect 42 -27 49 -23
rect 38 -28 46 -27
rect 38 -30 39 -28
rect 41 -30 46 -28
rect 38 -31 46 -30
<< ptie >>
rect -9 30 -3 32
rect -9 28 -7 30
rect -5 28 -3 30
rect -9 26 -3 28
rect 53 30 59 32
rect 53 28 55 30
rect 57 28 59 30
rect 53 26 59 28
rect -9 0 -3 2
rect -9 -2 -7 0
rect -5 -2 -3 0
rect -9 -4 -3 -2
<< ntie >>
rect -53 90 -47 92
rect -53 88 -51 90
rect -49 88 -47 90
rect -53 86 -47 88
rect -53 -60 -47 -58
rect -53 -62 -51 -60
rect -49 -62 -47 -60
rect -53 -64 -47 -62
<< nmos >>
rect -41 29 -39 49
rect -31 29 -29 49
rect -21 29 -19 49
rect -11 40 -9 49
rect 15 36 17 49
rect 22 36 24 49
rect 35 35 37 49
rect 59 38 61 46
rect 70 35 72 43
rect -41 -21 -39 -1
rect -31 -21 -29 -1
rect -21 -21 -19 -1
rect -11 -21 -9 -12
rect 13 -21 15 -8
rect 20 -21 22 -8
rect 33 -21 35 -7
<< pmos >>
rect -41 61 -39 81
rect -31 61 -29 89
rect -21 61 -19 89
rect -11 61 -9 89
rect 15 70 17 89
rect 25 70 27 89
rect 35 61 37 89
rect 61 61 63 89
rect 68 61 70 89
rect -41 -53 -39 -33
rect -31 -61 -29 -33
rect -21 -61 -19 -33
rect -11 -61 -9 -33
rect 13 -61 15 -42
rect 23 -61 25 -42
rect 33 -61 35 -33
<< polyct0 >>
rect 33 54 35 56
rect 31 -28 33 -26
<< polyct1 >>
rect 13 62 15 64
rect -39 54 -37 56
rect -31 54 -29 56
rect 23 54 25 56
rect 59 51 61 53
rect 69 54 71 56
rect -39 -28 -37 -26
rect -31 -28 -29 -26
rect 21 -28 23 -26
rect 11 -36 13 -34
<< ndifct0 >>
rect -47 38 -45 40
rect -47 31 -45 33
rect -26 38 -24 40
rect -26 31 -24 33
rect -6 42 -4 44
rect 10 38 12 40
rect 54 40 56 42
rect -47 -5 -45 -3
rect -47 -12 -45 -10
rect -26 -5 -24 -3
rect -26 -12 -24 -10
rect 8 -12 10 -10
rect -6 -16 -4 -14
<< ndifct1 >>
rect -36 45 -34 47
rect -36 38 -34 40
rect -16 45 -14 47
rect 40 45 42 47
rect 40 37 42 39
rect 65 37 67 39
rect 29 28 31 30
rect 76 28 78 30
rect -36 -12 -34 -10
rect -36 -19 -34 -17
rect 27 -2 29 0
rect -16 -19 -14 -17
rect 38 -11 40 -9
rect 38 -19 40 -17
<< ntiect1 >>
rect -51 88 -49 90
rect -51 -62 -49 -60
<< ptiect1 >>
rect -7 28 -5 30
rect 55 28 57 30
rect -7 -2 -5 0
<< pdifct0 >>
rect -46 77 -44 79
rect -46 70 -44 72
rect -26 85 -24 87
rect -26 77 -24 79
rect -16 70 -14 72
rect -6 85 -4 87
rect -6 78 -4 80
rect 10 85 12 87
rect 10 78 12 80
rect 20 79 22 81
rect 20 72 22 74
rect 30 85 32 87
rect 30 78 32 80
rect 54 85 56 87
rect 54 78 56 80
rect -46 -44 -44 -42
rect -46 -51 -44 -49
rect -26 -51 -24 -49
rect -26 -59 -24 -57
rect -16 -44 -14 -42
rect -6 -52 -4 -50
rect -6 -59 -4 -57
rect 8 -52 10 -50
rect 8 -59 10 -57
rect 18 -46 20 -44
rect 18 -53 20 -51
rect 28 -52 30 -50
rect 28 -59 30 -57
<< pdifct1 >>
rect -36 70 -34 72
rect -36 63 -34 65
rect -16 63 -14 65
rect 40 78 42 80
rect 40 71 42 73
rect 73 78 75 80
rect 73 71 75 73
rect -36 -37 -34 -35
rect -36 -44 -34 -42
rect -16 -37 -14 -35
rect 38 -45 40 -43
rect 38 -52 40 -50
<< alu0 >>
rect -48 79 -42 87
rect -48 77 -46 79
rect -44 77 -42 79
rect -48 72 -42 77
rect -27 85 -26 87
rect -24 85 -23 87
rect -27 79 -23 85
rect -27 77 -26 79
rect -24 77 -23 79
rect -8 85 -6 87
rect -4 85 -2 87
rect -8 80 -2 85
rect -8 78 -6 80
rect -4 78 -2 80
rect -8 77 -2 78
rect 8 85 10 87
rect 12 85 14 87
rect 8 80 14 85
rect 28 85 30 87
rect 32 85 34 87
rect 8 78 10 80
rect 12 78 14 80
rect 8 77 14 78
rect 18 81 24 82
rect 18 79 20 81
rect 22 79 24 81
rect -27 75 -23 77
rect 18 74 24 79
rect 28 80 34 85
rect 53 85 54 87
rect 56 85 57 87
rect 28 78 30 80
rect 32 78 34 80
rect 28 77 34 78
rect -48 70 -46 72
rect -44 70 -42 72
rect -48 69 -42 70
rect -17 72 -13 74
rect -17 70 -16 72
rect -14 70 -13 72
rect -17 66 -13 70
rect -17 65 -14 66
rect 18 72 20 74
rect 22 73 24 74
rect 53 80 57 85
rect 53 78 54 80
rect 56 78 57 80
rect 53 76 57 78
rect 22 72 32 73
rect 18 69 32 72
rect 28 65 32 69
rect 28 61 36 65
rect 32 56 36 61
rect 32 54 33 56
rect 35 54 36 56
rect 32 49 36 54
rect -49 40 -43 41
rect -49 38 -47 40
rect -45 38 -43 40
rect -49 33 -43 38
rect -7 44 -3 46
rect 24 45 36 49
rect -7 42 -6 44
rect -4 42 -3 44
rect -28 40 -22 41
rect -28 38 -26 40
rect -24 38 -22 40
rect -49 31 -47 33
rect -45 31 -43 33
rect -28 33 -22 38
rect -28 31 -26 33
rect -24 31 -22 33
rect -7 31 -3 42
rect 24 41 28 45
rect 39 42 40 49
rect 8 40 28 41
rect 8 38 10 40
rect 12 38 28 40
rect 8 37 28 38
rect 53 42 57 44
rect 53 40 54 42
rect 56 40 57 42
rect 53 31 57 40
rect -49 -5 -47 -3
rect -45 -5 -43 -3
rect -49 -10 -43 -5
rect -28 -5 -26 -3
rect -24 -5 -22 -3
rect -49 -12 -47 -10
rect -45 -12 -43 -10
rect -49 -13 -43 -12
rect -28 -10 -22 -5
rect -28 -12 -26 -10
rect -24 -12 -22 -10
rect -28 -13 -22 -12
rect -7 -14 -3 -3
rect 6 -10 26 -9
rect 6 -12 8 -10
rect 10 -12 26 -10
rect 6 -13 26 -12
rect -7 -16 -6 -14
rect -4 -16 -3 -14
rect -7 -18 -3 -16
rect 22 -17 26 -13
rect 22 -21 34 -17
rect 37 -21 38 -14
rect 30 -26 34 -21
rect 30 -28 31 -26
rect 33 -28 34 -26
rect 30 -33 34 -28
rect 26 -37 34 -33
rect -48 -42 -42 -41
rect -48 -44 -46 -42
rect -44 -44 -42 -42
rect -48 -49 -42 -44
rect -17 -38 -14 -37
rect -17 -42 -13 -38
rect -17 -44 -16 -42
rect -14 -44 -13 -42
rect -17 -46 -13 -44
rect 26 -41 30 -37
rect 16 -44 30 -41
rect 16 -46 18 -44
rect 20 -45 30 -44
rect 20 -46 22 -45
rect -48 -51 -46 -49
rect -44 -51 -42 -49
rect -48 -59 -42 -51
rect -27 -49 -23 -47
rect -27 -51 -26 -49
rect -24 -51 -23 -49
rect -27 -57 -23 -51
rect -27 -59 -26 -57
rect -24 -59 -23 -57
rect -8 -50 -2 -49
rect -8 -52 -6 -50
rect -4 -52 -2 -50
rect -8 -57 -2 -52
rect -8 -59 -6 -57
rect -4 -59 -2 -57
rect 6 -50 12 -49
rect 6 -52 8 -50
rect 10 -52 12 -50
rect 6 -57 12 -52
rect 16 -51 22 -46
rect 16 -53 18 -51
rect 20 -53 22 -51
rect 16 -54 22 -53
rect 26 -50 32 -49
rect 26 -52 28 -50
rect 30 -52 32 -50
rect 6 -59 8 -57
rect 10 -59 12 -57
rect 26 -57 32 -52
rect 26 -59 28 -57
rect 30 -59 32 -57
<< via1 >>
rect -59 55 -57 57
rect 17 45 19 47
rect 49 51 51 53
rect -49 -28 -47 -26
rect 2 -28 4 -26
rect 39 -30 41 -28
<< via2 >>
rect 49 51 51 53
rect 17 45 19 47
rect -49 -28 -47 -26
rect 39 -30 41 -28
<< via3 >>
rect 49 51 51 53
rect 39 -30 41 -28
<< labels >>
rlabel alu1 -45 55 -45 55 1 A
rlabel alu1 -12 53 -12 53 1 -A
rlabel alu1 10 64 10 64 1 -A
rlabel alu1 19 54 19 54 1 B
rlabel alu0 33 59 33 59 1 and_a_b_node
rlabel alu1 -44 -26 -44 -26 1 B
rlabel alu1 -13 -25 -13 -25 1 -B
rlabel alu1 8 -39 8 -39 1 -B
rlabel alu1 16 -24 16 -24 1 A
rlabel alu0 31 -23 31 -23 1 and_a_b_node2
rlabel alu1 78 53 78 53 3 fout_1bit
rlabel alu1 40 -26 40 -26 1 GT_1bit
rlabel alu1 40 56 44 60 1 LT_1bit
rlabel nwell -57 87 82 95 1 vdd
rlabel alu1 -10 26 -10 27 1 vss
<< end >>
