magic
tech scmos
timestamp 1635784308
<< nwell >>
rect -8 -4 7 13
<< polysilicon >>
rect -1 4 1 6
rect -1 -5 1 -2
rect 0 -9 1 -5
rect -1 -12 1 -9
rect -1 -17 1 -15
<< ndiffusion >>
rect -2 -15 -1 -12
rect 1 -15 3 -12
<< pdiffusion >>
rect -4 3 -1 4
rect -2 -1 -1 3
rect -4 -2 -1 -1
rect 1 3 4 4
rect 1 -1 2 3
rect 1 -2 4 -1
<< metal1 >>
rect -2 9 2 12
rect -6 3 -3 9
rect 3 -5 6 -1
rect -7 -9 -4 -5
rect 3 -8 9 -5
rect 3 -12 6 -8
rect -5 -19 -2 -16
rect -5 -20 6 -19
rect -1 -22 3 -20
<< ntransistor >>
rect -1 -15 1 -12
<< ptransistor >>
rect -1 -2 1 4
<< polycontact >>
rect -4 -9 0 -5
<< ndcontact >>
rect -6 -16 -2 -12
rect 3 -16 7 -12
<< pdcontact >>
rect -6 -1 -2 3
rect 2 -1 6 3
<< psubstratepcontact >>
rect -5 -24 -1 -20
rect 3 -24 7 -20
<< nsubstratencontact >>
rect -6 9 -2 13
rect 2 9 6 13
<< labels >>
rlabel metal1 1 -21 1 -21 1 gnd
rlabel metal1 6 -7 6 -7 1 out
rlabel metal1 -5 -7 -5 -7 1 in
rlabel metal1 0 11 0 11 1 V_DD
<< end >>
