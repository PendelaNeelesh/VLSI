magic
tech scmos
timestamp 1635821822
<< nwell >>
rect -17 18 22 34
<< polysilicon >>
rect 0 26 2 28
rect 10 26 12 28
rect 0 18 2 20
rect -8 17 2 18
rect -7 16 2 17
rect 10 17 12 20
rect -7 13 -6 16
rect 10 14 11 17
rect -8 10 -6 13
rect -2 13 11 14
rect -2 12 12 13
rect -2 10 0 12
rect -8 5 -6 7
rect -2 5 0 7
<< ndiffusion >>
rect -10 7 -8 10
rect -6 7 -2 10
rect 0 7 2 10
<< pdiffusion >>
rect -4 25 0 26
rect -2 20 0 25
rect 2 25 10 26
rect 2 20 4 25
rect 8 20 10 25
rect 12 25 16 26
rect 12 20 14 25
<< metal1 >>
rect -17 30 -14 34
rect -10 30 -6 34
rect -2 30 2 34
rect 6 30 11 34
rect 15 30 22 34
rect -6 25 -2 30
rect 15 25 19 30
rect 3 20 4 22
rect 18 20 19 25
rect -14 13 -11 17
rect 3 10 7 20
rect 15 13 19 17
rect 6 6 19 10
rect -14 1 -10 6
rect -17 -2 -14 1
rect -10 -2 -6 1
rect -2 -2 2 1
rect 6 -2 11 1
rect 15 -2 22 1
<< ntransistor >>
rect -8 7 -6 10
rect -2 7 0 10
<< ptransistor >>
rect 0 20 2 26
rect 10 20 12 26
<< polycontact >>
rect -11 13 -7 17
rect 11 13 15 17
<< ndcontact >>
rect -14 6 -10 10
rect 2 6 6 10
<< pdcontact >>
rect -6 20 -2 25
rect 4 20 8 25
rect 14 20 18 25
<< psubstratepcontact >>
rect -14 -3 -10 1
rect -6 -3 -2 1
rect 2 -3 6 1
rect 11 -3 15 1
<< nsubstratencontact >>
rect -14 30 -10 35
rect -6 30 -2 35
rect 2 30 6 35
rect 11 30 15 35
<< labels >>
rlabel metal1 0 32 0 32 5 V_DD
rlabel metal1 0 -1 0 -1 1 gnd
rlabel metal1 -13 15 -13 15 3 A
rlabel metal1 17 15 17 15 7 B
rlabel metal1 17 8 17 8 7 out
rlabel ndiffusion -4 9 -4 9 1 pdn_a_b
<< end >>
