magic
tech scmos
timestamp 1636124730
<< ab >>
rect -11 192 29 264
rect 33 192 73 264
rect 83 192 123 264
rect 133 192 173 264
rect 183 192 231 264
rect -7 91 49 163
rect 55 127 95 163
rect 99 127 131 163
rect 55 123 93 127
rect 55 91 95 123
rect 99 122 101 123
rect 105 122 131 127
rect 99 91 131 122
rect 133 91 173 163
rect 177 91 233 163
rect -7 1 49 73
rect 53 1 93 73
rect 95 42 127 73
rect 95 37 121 42
rect 125 41 127 42
rect 131 41 171 73
rect 133 37 171 41
rect 95 1 127 37
rect 131 1 171 37
rect 177 1 233 73
<< nwell >>
rect -16 187 236 232
rect -12 123 238 168
rect -12 6 238 41
rect 95 -4 238 6
<< pwell >>
rect -16 232 236 269
rect -12 91 238 123
rect -12 41 238 73
<< poly >>
rect -2 252 0 257
rect 8 251 10 256
rect 18 249 20 253
rect 42 252 44 257
rect -2 235 0 238
rect 8 235 10 243
rect 18 235 20 241
rect 55 251 57 256
rect 62 251 64 256
rect 92 252 94 257
rect 102 251 104 256
rect 208 258 210 262
rect 218 258 220 262
rect 112 249 114 253
rect 142 251 144 256
rect 149 251 151 256
rect 162 252 164 257
rect 42 235 44 238
rect 55 235 57 238
rect -2 233 4 235
rect -2 231 0 233
rect 2 231 4 233
rect -2 229 4 231
rect 8 233 14 235
rect 8 231 10 233
rect 12 231 14 233
rect 8 229 14 231
rect 18 233 27 235
rect 18 231 23 233
rect 25 231 27 233
rect 18 229 27 231
rect 42 233 48 235
rect 42 231 44 233
rect 46 231 48 233
rect 42 229 48 231
rect 52 233 58 235
rect 52 231 54 233
rect 56 231 58 233
rect 52 229 58 231
rect -2 226 0 229
rect 11 226 13 229
rect 18 226 20 229
rect 42 226 44 229
rect -2 194 0 198
rect 52 217 54 229
rect 62 227 64 238
rect 92 235 94 238
rect 102 235 104 243
rect 112 235 114 241
rect 192 241 198 243
rect 192 239 194 241
rect 196 239 198 241
rect 92 233 98 235
rect 92 231 94 233
rect 96 231 98 233
rect 92 229 98 231
rect 102 233 108 235
rect 102 231 104 233
rect 106 231 108 233
rect 102 229 108 231
rect 112 233 121 235
rect 112 231 117 233
rect 119 231 121 233
rect 112 229 121 231
rect 62 225 68 227
rect 92 226 94 229
rect 105 226 107 229
rect 112 226 114 229
rect 142 227 144 238
rect 149 235 151 238
rect 162 235 164 238
rect 192 237 198 239
rect 148 233 154 235
rect 148 231 150 233
rect 152 231 154 233
rect 148 229 154 231
rect 158 233 164 235
rect 158 231 160 233
rect 162 231 164 233
rect 158 229 164 231
rect 62 223 64 225
rect 66 223 68 225
rect 62 221 68 223
rect 62 217 64 221
rect 11 194 13 198
rect 18 194 20 198
rect 42 194 44 198
rect 52 194 54 198
rect 62 194 64 198
rect 92 194 94 198
rect 138 225 144 227
rect 138 223 140 225
rect 142 223 144 225
rect 138 221 144 223
rect 142 217 144 221
rect 152 217 154 229
rect 162 226 164 229
rect 196 225 198 237
rect 208 235 210 243
rect 218 240 220 243
rect 203 233 210 235
rect 214 238 220 240
rect 214 236 216 238
rect 218 237 220 238
rect 218 236 222 237
rect 214 234 222 236
rect 203 231 205 233
rect 207 231 210 233
rect 203 230 210 231
rect 203 228 215 230
rect 203 225 205 228
rect 213 225 215 228
rect 220 225 222 234
rect 105 194 107 198
rect 112 194 114 198
rect 142 194 144 198
rect 152 194 154 198
rect 162 194 164 198
rect 196 194 198 198
rect 203 194 205 198
rect 213 194 215 198
rect 220 194 222 198
rect 18 157 20 161
rect 28 157 30 161
rect 38 157 40 161
rect 64 157 66 161
rect 74 157 76 161
rect 84 157 86 161
rect 110 157 112 161
rect 117 157 119 161
rect 142 157 144 161
rect 152 157 154 161
rect 162 157 164 161
rect 186 157 188 161
rect 196 157 198 161
rect 206 157 208 161
rect 8 149 10 153
rect 64 134 66 138
rect 60 132 66 134
rect 60 130 62 132
rect 64 130 66 132
rect 8 126 10 129
rect 18 126 20 129
rect 28 126 30 129
rect 38 126 40 129
rect 60 128 66 130
rect 8 124 40 126
rect 8 122 10 124
rect 12 122 18 124
rect 20 122 22 124
rect 8 120 22 122
rect 8 117 10 120
rect 18 117 20 120
rect 28 117 30 124
rect 38 117 40 124
rect 64 117 66 128
rect 74 126 76 138
rect 84 126 86 129
rect 70 124 76 126
rect 70 122 72 124
rect 74 122 76 124
rect 70 120 76 122
rect 80 124 86 126
rect 80 122 82 124
rect 84 122 86 124
rect 110 123 112 129
rect 117 126 119 129
rect 142 126 144 129
rect 152 126 154 138
rect 162 134 164 138
rect 162 132 168 134
rect 162 130 164 132
rect 166 130 168 132
rect 162 128 168 130
rect 216 149 218 153
rect 80 120 86 122
rect 71 117 73 120
rect 84 117 86 120
rect 106 121 112 123
rect 106 119 108 121
rect 110 119 112 121
rect 116 124 122 126
rect 116 122 118 124
rect 120 122 122 124
rect 116 120 122 122
rect 142 124 148 126
rect 142 122 144 124
rect 146 122 148 124
rect 142 120 148 122
rect 152 124 158 126
rect 152 122 154 124
rect 156 122 158 124
rect 152 120 158 122
rect 106 117 112 119
rect 38 103 40 108
rect 64 99 66 104
rect 71 99 73 104
rect 108 114 110 117
rect 119 111 121 120
rect 142 117 144 120
rect 155 117 157 120
rect 162 117 164 128
rect 186 126 188 129
rect 196 126 198 129
rect 206 126 208 129
rect 216 126 218 129
rect 186 124 218 126
rect 186 117 188 124
rect 196 117 198 124
rect 204 122 206 124
rect 208 122 214 124
rect 216 122 218 124
rect 204 120 218 122
rect 206 117 208 120
rect 216 117 218 120
rect 8 93 10 97
rect 18 93 20 97
rect 28 93 30 97
rect 84 98 86 103
rect 108 102 110 106
rect 119 98 121 103
rect 142 98 144 103
rect 155 99 157 104
rect 162 99 164 104
rect 186 103 188 108
rect 196 93 198 97
rect 206 93 208 97
rect 216 93 218 97
rect 8 67 10 71
rect 18 67 20 71
rect 28 67 30 71
rect 38 56 40 61
rect 62 60 64 65
rect 69 60 71 65
rect 82 61 84 66
rect 105 61 107 66
rect 116 58 118 62
rect 140 61 142 66
rect 196 67 198 71
rect 206 67 208 71
rect 216 67 218 71
rect 8 44 10 47
rect 18 44 20 47
rect 8 42 22 44
rect 8 40 10 42
rect 12 40 18 42
rect 20 40 22 42
rect 28 40 30 47
rect 38 40 40 47
rect 8 38 40 40
rect 8 35 10 38
rect 18 35 20 38
rect 28 35 30 38
rect 38 35 40 38
rect 62 36 64 47
rect 69 44 71 47
rect 82 44 84 47
rect 105 44 107 53
rect 116 47 118 50
rect 153 60 155 65
rect 160 60 162 65
rect 186 56 188 61
rect 114 45 120 47
rect 68 42 74 44
rect 68 40 70 42
rect 72 40 74 42
rect 68 38 74 40
rect 78 42 84 44
rect 78 40 80 42
rect 82 40 84 42
rect 78 38 84 40
rect 104 42 110 44
rect 104 40 106 42
rect 108 40 110 42
rect 104 38 110 40
rect 114 43 116 45
rect 118 43 120 45
rect 114 41 120 43
rect 140 44 142 47
rect 153 44 155 47
rect 140 42 146 44
rect 8 11 10 15
rect 58 34 64 36
rect 58 32 60 34
rect 62 32 64 34
rect 58 30 64 32
rect 62 26 64 30
rect 72 26 74 38
rect 82 35 84 38
rect 107 35 109 38
rect 114 35 116 41
rect 140 40 142 42
rect 144 40 146 42
rect 140 38 146 40
rect 150 42 156 44
rect 150 40 152 42
rect 154 40 156 42
rect 150 38 156 40
rect 140 35 142 38
rect 150 26 152 38
rect 160 36 162 47
rect 186 40 188 47
rect 196 40 198 47
rect 206 44 208 47
rect 216 44 218 47
rect 204 42 218 44
rect 204 40 206 42
rect 208 40 214 42
rect 216 40 218 42
rect 186 38 218 40
rect 160 34 166 36
rect 186 35 188 38
rect 196 35 198 38
rect 206 35 208 38
rect 216 35 218 38
rect 160 32 162 34
rect 164 32 166 34
rect 160 30 166 32
rect 160 26 162 30
rect 216 11 218 15
rect 18 3 20 7
rect 28 3 30 7
rect 38 3 40 7
rect 62 3 64 7
rect 72 3 74 7
rect 82 3 84 7
rect 107 3 109 7
rect 114 3 116 7
rect 140 3 142 7
rect 150 3 152 7
rect 160 3 162 7
rect 186 3 188 7
rect 196 3 198 7
rect 206 3 208 7
<< ndif >>
rect 46 259 53 261
rect 46 257 48 259
rect 50 257 53 259
rect -9 249 -2 252
rect -9 247 -7 249
rect -5 247 -2 249
rect -9 242 -2 247
rect -9 240 -7 242
rect -5 240 -2 242
rect -9 238 -2 240
rect 0 251 5 252
rect 0 249 8 251
rect 0 247 3 249
rect 5 247 8 249
rect 0 243 8 247
rect 10 249 15 251
rect 46 252 53 257
rect 35 250 42 252
rect 10 247 18 249
rect 10 245 13 247
rect 15 245 18 247
rect 10 243 18 245
rect 0 238 5 243
rect 13 241 18 243
rect 20 247 27 249
rect 20 245 23 247
rect 25 245 27 247
rect 20 241 27 245
rect 35 248 37 250
rect 39 248 42 250
rect 35 242 42 248
rect 35 240 37 242
rect 39 240 42 242
rect 35 238 42 240
rect 44 251 53 252
rect 44 238 55 251
rect 57 238 62 251
rect 64 249 71 251
rect 64 247 67 249
rect 69 247 71 249
rect 64 245 71 247
rect 85 249 92 252
rect 85 247 87 249
rect 89 247 92 249
rect 64 238 69 245
rect 85 242 92 247
rect 85 240 87 242
rect 89 240 92 242
rect 85 238 92 240
rect 94 251 99 252
rect 153 259 160 261
rect 153 257 156 259
rect 158 257 160 259
rect 94 249 102 251
rect 94 247 97 249
rect 99 247 102 249
rect 94 243 102 247
rect 104 249 109 251
rect 153 252 160 257
rect 153 251 162 252
rect 135 249 142 251
rect 104 247 112 249
rect 104 245 107 247
rect 109 245 112 247
rect 104 243 112 245
rect 94 238 99 243
rect 107 241 112 243
rect 114 247 121 249
rect 114 245 117 247
rect 119 245 121 247
rect 135 247 137 249
rect 139 247 142 249
rect 135 245 142 247
rect 114 241 121 245
rect 137 238 142 245
rect 144 238 149 251
rect 151 238 162 251
rect 164 250 171 252
rect 164 248 167 250
rect 169 248 171 250
rect 164 242 171 248
rect 200 256 208 258
rect 200 254 203 256
rect 205 254 208 256
rect 200 249 208 254
rect 200 247 203 249
rect 205 247 208 249
rect 200 243 208 247
rect 210 249 218 258
rect 210 247 213 249
rect 215 247 218 249
rect 210 243 218 247
rect 220 256 228 258
rect 220 254 223 256
rect 225 254 228 256
rect 220 243 228 254
rect 164 240 167 242
rect 169 240 171 242
rect 164 238 171 240
rect 0 108 8 117
rect 0 106 2 108
rect 4 106 8 108
rect 0 101 8 106
rect 0 99 2 101
rect 4 99 8 101
rect 0 97 8 99
rect 10 115 18 117
rect 10 113 13 115
rect 15 113 18 115
rect 10 108 18 113
rect 10 106 13 108
rect 15 106 18 108
rect 10 97 18 106
rect 20 108 28 117
rect 20 106 23 108
rect 25 106 28 108
rect 20 101 28 106
rect 20 99 23 101
rect 25 99 28 101
rect 20 97 28 99
rect 30 115 38 117
rect 30 113 33 115
rect 35 113 38 115
rect 30 108 38 113
rect 40 112 47 117
rect 40 110 43 112
rect 45 110 47 112
rect 59 110 64 117
rect 40 108 47 110
rect 57 108 64 110
rect 30 97 35 108
rect 57 106 59 108
rect 61 106 64 108
rect 57 104 64 106
rect 66 104 71 117
rect 73 104 84 117
rect 75 103 84 104
rect 86 115 93 117
rect 86 113 89 115
rect 91 113 93 115
rect 86 107 93 113
rect 86 105 89 107
rect 91 105 93 107
rect 101 110 108 114
rect 101 108 103 110
rect 105 108 108 110
rect 101 106 108 108
rect 110 111 115 114
rect 135 115 142 117
rect 135 113 137 115
rect 139 113 142 115
rect 110 107 119 111
rect 110 106 114 107
rect 86 103 93 105
rect 75 98 82 103
rect 112 105 114 106
rect 116 105 119 107
rect 112 103 119 105
rect 121 103 129 111
rect 135 107 142 113
rect 135 105 137 107
rect 139 105 142 107
rect 135 103 142 105
rect 144 104 155 117
rect 157 104 162 117
rect 164 110 169 117
rect 179 112 186 117
rect 179 110 181 112
rect 183 110 186 112
rect 164 108 171 110
rect 179 108 186 110
rect 188 115 196 117
rect 188 113 191 115
rect 193 113 196 115
rect 188 108 196 113
rect 164 106 167 108
rect 169 106 171 108
rect 164 104 171 106
rect 144 103 153 104
rect 123 98 129 103
rect 146 98 153 103
rect 75 96 78 98
rect 80 96 82 98
rect 75 94 82 96
rect 123 96 125 98
rect 127 96 129 98
rect 123 94 129 96
rect 146 96 148 98
rect 150 96 153 98
rect 146 94 153 96
rect 191 97 196 108
rect 198 108 206 117
rect 198 106 201 108
rect 203 106 206 108
rect 198 101 206 106
rect 198 99 201 101
rect 203 99 206 101
rect 198 97 206 99
rect 208 115 216 117
rect 208 113 211 115
rect 213 113 216 115
rect 208 108 216 113
rect 208 106 211 108
rect 213 106 216 108
rect 208 97 216 106
rect 218 108 226 117
rect 218 106 222 108
rect 224 106 226 108
rect 218 101 226 106
rect 218 99 222 101
rect 224 99 226 101
rect 218 97 226 99
rect 0 65 8 67
rect 0 63 2 65
rect 4 63 8 65
rect 0 58 8 63
rect 0 56 2 58
rect 4 56 8 58
rect 0 47 8 56
rect 10 58 18 67
rect 10 56 13 58
rect 15 56 18 58
rect 10 51 18 56
rect 10 49 13 51
rect 15 49 18 51
rect 10 47 18 49
rect 20 65 28 67
rect 20 63 23 65
rect 25 63 28 65
rect 20 58 28 63
rect 20 56 23 58
rect 25 56 28 58
rect 20 47 28 56
rect 30 56 35 67
rect 73 68 80 70
rect 73 66 76 68
rect 78 66 80 68
rect 97 68 103 70
rect 97 66 99 68
rect 101 66 103 68
rect 144 68 151 70
rect 144 66 146 68
rect 148 66 151 68
rect 73 61 80 66
rect 97 61 103 66
rect 73 60 82 61
rect 55 58 62 60
rect 55 56 57 58
rect 59 56 62 58
rect 30 51 38 56
rect 30 49 33 51
rect 35 49 38 51
rect 30 47 38 49
rect 40 54 47 56
rect 55 54 62 56
rect 40 52 43 54
rect 45 52 47 54
rect 40 47 47 52
rect 57 47 62 54
rect 64 47 69 60
rect 71 47 82 60
rect 84 59 91 61
rect 84 57 87 59
rect 89 57 91 59
rect 84 51 91 57
rect 97 53 105 61
rect 107 59 114 61
rect 107 57 110 59
rect 112 58 114 59
rect 144 61 151 66
rect 133 59 140 61
rect 112 57 116 58
rect 107 53 116 57
rect 84 49 87 51
rect 89 49 91 51
rect 84 47 91 49
rect 111 50 116 53
rect 118 56 125 58
rect 118 54 121 56
rect 123 54 125 56
rect 118 50 125 54
rect 133 57 135 59
rect 137 57 140 59
rect 133 51 140 57
rect 133 49 135 51
rect 137 49 140 51
rect 133 47 140 49
rect 142 60 151 61
rect 142 47 153 60
rect 155 47 160 60
rect 162 58 169 60
rect 162 56 165 58
rect 167 56 169 58
rect 191 56 196 67
rect 162 54 169 56
rect 179 54 186 56
rect 162 47 167 54
rect 179 52 181 54
rect 183 52 186 54
rect 179 47 186 52
rect 188 51 196 56
rect 188 49 191 51
rect 193 49 196 51
rect 188 47 196 49
rect 198 65 206 67
rect 198 63 201 65
rect 203 63 206 65
rect 198 58 206 63
rect 198 56 201 58
rect 203 56 206 58
rect 198 47 206 56
rect 208 58 216 67
rect 208 56 211 58
rect 213 56 216 58
rect 208 51 216 56
rect 208 49 211 51
rect 213 49 216 51
rect 208 47 216 49
rect 218 65 226 67
rect 218 63 222 65
rect 224 63 226 65
rect 218 58 226 63
rect 218 56 222 58
rect 224 56 226 58
rect 218 47 226 56
<< pdif >>
rect -7 217 -2 226
rect -9 215 -2 217
rect -9 213 -7 215
rect -5 213 -2 215
rect -9 208 -2 213
rect -9 206 -7 208
rect -5 206 -2 208
rect -9 204 -2 206
rect -7 198 -2 204
rect 0 199 11 226
rect 0 198 4 199
rect 2 197 4 198
rect 6 198 11 199
rect 13 198 18 226
rect 20 210 25 226
rect 37 218 42 226
rect 35 216 42 218
rect 35 214 37 216
rect 39 214 42 216
rect 20 208 27 210
rect 20 206 23 208
rect 25 206 27 208
rect 20 204 27 206
rect 35 209 42 214
rect 35 207 37 209
rect 39 207 42 209
rect 35 205 42 207
rect 20 198 25 204
rect 37 198 42 205
rect 44 217 50 226
rect 87 217 92 226
rect 44 209 52 217
rect 44 207 47 209
rect 49 207 52 209
rect 44 202 52 207
rect 44 200 47 202
rect 49 200 52 202
rect 44 198 52 200
rect 54 215 62 217
rect 54 213 57 215
rect 59 213 62 215
rect 54 208 62 213
rect 54 206 57 208
rect 59 206 62 208
rect 54 198 62 206
rect 64 209 71 217
rect 64 207 67 209
rect 69 207 71 209
rect 64 202 71 207
rect 85 215 92 217
rect 85 213 87 215
rect 89 213 92 215
rect 85 208 92 213
rect 85 206 87 208
rect 89 206 92 208
rect 85 204 92 206
rect 64 200 67 202
rect 69 200 71 202
rect 64 198 71 200
rect 87 198 92 204
rect 94 199 105 226
rect 94 198 98 199
rect 6 197 9 198
rect 2 195 9 197
rect 96 197 98 198
rect 100 198 105 199
rect 107 198 112 226
rect 114 210 119 226
rect 156 217 162 226
rect 114 208 121 210
rect 114 206 117 208
rect 119 206 121 208
rect 114 204 121 206
rect 135 209 142 217
rect 135 207 137 209
rect 139 207 142 209
rect 114 198 119 204
rect 135 202 142 207
rect 135 200 137 202
rect 139 200 142 202
rect 135 198 142 200
rect 144 215 152 217
rect 144 213 147 215
rect 149 213 152 215
rect 144 208 152 213
rect 144 206 147 208
rect 149 206 152 208
rect 144 198 152 206
rect 154 209 162 217
rect 154 207 157 209
rect 159 207 162 209
rect 154 202 162 207
rect 154 200 157 202
rect 159 200 162 202
rect 154 198 162 200
rect 164 218 169 226
rect 164 216 171 218
rect 164 214 167 216
rect 169 214 171 216
rect 164 209 171 214
rect 164 207 167 209
rect 169 207 171 209
rect 164 205 171 207
rect 189 209 196 225
rect 189 207 191 209
rect 193 207 196 209
rect 164 198 169 205
rect 189 202 196 207
rect 189 200 191 202
rect 193 200 196 202
rect 189 198 196 200
rect 198 198 203 225
rect 205 223 213 225
rect 205 221 208 223
rect 210 221 213 223
rect 205 216 213 221
rect 205 214 208 216
rect 210 214 213 216
rect 205 198 213 214
rect 215 198 220 225
rect 222 209 229 225
rect 222 207 225 209
rect 227 207 229 209
rect 222 202 229 207
rect 222 200 225 202
rect 227 200 229 202
rect 222 198 229 200
rect 100 197 103 198
rect 96 195 103 197
rect 13 149 18 157
rect 1 147 8 149
rect 1 145 3 147
rect 5 145 8 147
rect 1 140 8 145
rect 1 138 3 140
rect 5 138 8 140
rect 1 129 8 138
rect 10 140 18 149
rect 10 138 13 140
rect 15 138 18 140
rect 10 133 18 138
rect 10 131 13 133
rect 15 131 18 133
rect 10 129 18 131
rect 20 155 28 157
rect 20 153 23 155
rect 25 153 28 155
rect 20 147 28 153
rect 20 145 23 147
rect 25 145 28 147
rect 20 129 28 145
rect 30 140 38 157
rect 30 138 33 140
rect 35 138 38 140
rect 30 133 38 138
rect 30 131 33 133
rect 35 131 38 133
rect 30 129 38 131
rect 40 155 47 157
rect 40 153 43 155
rect 45 153 47 155
rect 40 148 47 153
rect 40 146 43 148
rect 45 146 47 148
rect 40 129 47 146
rect 57 155 64 157
rect 57 153 59 155
rect 61 153 64 155
rect 57 148 64 153
rect 57 146 59 148
rect 61 146 64 148
rect 57 138 64 146
rect 66 149 74 157
rect 66 147 69 149
rect 71 147 74 149
rect 66 142 74 147
rect 66 140 69 142
rect 71 140 74 142
rect 66 138 74 140
rect 76 155 84 157
rect 76 153 79 155
rect 81 153 84 155
rect 76 148 84 153
rect 76 146 79 148
rect 81 146 84 148
rect 76 138 84 146
rect 78 129 84 138
rect 86 150 91 157
rect 101 155 110 157
rect 101 153 103 155
rect 105 153 110 155
rect 86 148 93 150
rect 86 146 89 148
rect 91 146 93 148
rect 86 141 93 146
rect 86 139 89 141
rect 91 139 93 141
rect 86 137 93 139
rect 101 148 110 153
rect 101 146 103 148
rect 105 146 110 148
rect 86 129 91 137
rect 101 129 110 146
rect 112 129 117 157
rect 119 150 124 157
rect 137 150 142 157
rect 119 148 126 150
rect 119 146 122 148
rect 124 146 126 148
rect 119 141 126 146
rect 119 139 122 141
rect 124 139 126 141
rect 119 137 126 139
rect 135 148 142 150
rect 135 146 137 148
rect 139 146 142 148
rect 135 141 142 146
rect 135 139 137 141
rect 139 139 142 141
rect 135 137 142 139
rect 119 129 124 137
rect 137 129 142 137
rect 144 155 152 157
rect 144 153 147 155
rect 149 153 152 155
rect 144 148 152 153
rect 144 146 147 148
rect 149 146 152 148
rect 144 138 152 146
rect 154 149 162 157
rect 154 147 157 149
rect 159 147 162 149
rect 154 142 162 147
rect 154 140 157 142
rect 159 140 162 142
rect 154 138 162 140
rect 164 155 171 157
rect 164 153 167 155
rect 169 153 171 155
rect 164 148 171 153
rect 164 146 167 148
rect 169 146 171 148
rect 164 138 171 146
rect 179 155 186 157
rect 179 153 181 155
rect 183 153 186 155
rect 179 148 186 153
rect 179 146 181 148
rect 183 146 186 148
rect 144 129 150 138
rect 179 129 186 146
rect 188 140 196 157
rect 188 138 191 140
rect 193 138 196 140
rect 188 133 196 138
rect 188 131 191 133
rect 193 131 196 133
rect 188 129 196 131
rect 198 155 206 157
rect 198 153 201 155
rect 203 153 206 155
rect 198 147 206 153
rect 198 145 201 147
rect 203 145 206 147
rect 198 129 206 145
rect 208 149 213 157
rect 208 140 216 149
rect 208 138 211 140
rect 213 138 216 140
rect 208 133 216 138
rect 208 131 211 133
rect 213 131 216 133
rect 208 129 216 131
rect 218 147 225 149
rect 218 145 221 147
rect 223 145 225 147
rect 218 140 225 145
rect 218 138 221 140
rect 223 138 225 140
rect 218 129 225 138
rect 1 26 8 35
rect 1 24 3 26
rect 5 24 8 26
rect 1 19 8 24
rect 1 17 3 19
rect 5 17 8 19
rect 1 15 8 17
rect 10 33 18 35
rect 10 31 13 33
rect 15 31 18 33
rect 10 26 18 31
rect 10 24 13 26
rect 15 24 18 26
rect 10 15 18 24
rect 13 7 18 15
rect 20 19 28 35
rect 20 17 23 19
rect 25 17 28 19
rect 20 11 28 17
rect 20 9 23 11
rect 25 9 28 11
rect 20 7 28 9
rect 30 33 38 35
rect 30 31 33 33
rect 35 31 38 33
rect 30 26 38 31
rect 30 24 33 26
rect 35 24 38 26
rect 30 7 38 24
rect 40 18 47 35
rect 76 26 82 35
rect 40 16 43 18
rect 45 16 47 18
rect 40 11 47 16
rect 40 9 43 11
rect 45 9 47 11
rect 40 7 47 9
rect 55 18 62 26
rect 55 16 57 18
rect 59 16 62 18
rect 55 11 62 16
rect 55 9 57 11
rect 59 9 62 11
rect 55 7 62 9
rect 64 24 72 26
rect 64 22 67 24
rect 69 22 72 24
rect 64 17 72 22
rect 64 15 67 17
rect 69 15 72 17
rect 64 7 72 15
rect 74 18 82 26
rect 74 16 77 18
rect 79 16 82 18
rect 74 11 82 16
rect 74 9 77 11
rect 79 9 82 11
rect 74 7 82 9
rect 84 27 89 35
rect 102 27 107 35
rect 84 25 91 27
rect 84 23 87 25
rect 89 23 91 25
rect 84 18 91 23
rect 84 16 87 18
rect 89 16 91 18
rect 84 14 91 16
rect 100 25 107 27
rect 100 23 102 25
rect 104 23 107 25
rect 100 18 107 23
rect 100 16 102 18
rect 104 16 107 18
rect 100 14 107 16
rect 84 7 89 14
rect 102 7 107 14
rect 109 7 114 35
rect 116 18 125 35
rect 135 27 140 35
rect 116 16 121 18
rect 123 16 125 18
rect 116 11 125 16
rect 133 25 140 27
rect 133 23 135 25
rect 137 23 140 25
rect 133 18 140 23
rect 133 16 135 18
rect 137 16 140 18
rect 133 14 140 16
rect 116 9 121 11
rect 123 9 125 11
rect 116 7 125 9
rect 135 7 140 14
rect 142 26 148 35
rect 142 18 150 26
rect 142 16 145 18
rect 147 16 150 18
rect 142 11 150 16
rect 142 9 145 11
rect 147 9 150 11
rect 142 7 150 9
rect 152 24 160 26
rect 152 22 155 24
rect 157 22 160 24
rect 152 17 160 22
rect 152 15 155 17
rect 157 15 160 17
rect 152 7 160 15
rect 162 18 169 26
rect 162 16 165 18
rect 167 16 169 18
rect 162 11 169 16
rect 162 9 165 11
rect 167 9 169 11
rect 162 7 169 9
rect 179 18 186 35
rect 179 16 181 18
rect 183 16 186 18
rect 179 11 186 16
rect 179 9 181 11
rect 183 9 186 11
rect 179 7 186 9
rect 188 33 196 35
rect 188 31 191 33
rect 193 31 196 33
rect 188 26 196 31
rect 188 24 191 26
rect 193 24 196 26
rect 188 7 196 24
rect 198 19 206 35
rect 198 17 201 19
rect 203 17 206 19
rect 198 11 206 17
rect 198 9 201 11
rect 203 9 206 11
rect 198 7 206 9
rect 208 33 216 35
rect 208 31 211 33
rect 213 31 216 33
rect 208 26 216 31
rect 208 24 211 26
rect 213 24 216 26
rect 208 15 216 24
rect 218 26 225 35
rect 218 24 221 26
rect 223 24 225 26
rect 218 19 225 24
rect 218 17 221 19
rect 223 17 225 19
rect 218 15 225 17
rect 208 7 213 15
<< alu1 >>
rect 233 264 255 265
rect -13 259 255 264
rect -13 257 20 259
rect 22 257 48 259
rect 50 257 114 259
rect 116 257 156 259
rect 158 257 188 259
rect 190 257 255 259
rect -13 256 255 257
rect -9 249 -4 251
rect -9 247 -7 249
rect -5 247 -4 249
rect -9 242 -4 247
rect 35 250 47 251
rect 35 248 37 250
rect 39 248 47 250
rect 35 245 47 248
rect 85 249 90 251
rect 85 247 87 249
rect 89 247 90 249
rect 85 246 90 247
rect -9 240 -7 242
rect -5 240 -4 242
rect -9 238 -4 240
rect 35 242 39 245
rect 35 240 37 242
rect -9 234 -5 238
rect -9 232 -8 234
rect -6 232 -5 234
rect -9 215 -5 232
rect 7 233 19 235
rect 7 231 10 233
rect 12 231 19 233
rect 7 229 19 231
rect 7 227 11 229
rect 7 224 8 227
rect 10 224 11 227
rect 7 221 11 224
rect 23 233 27 235
rect 25 231 27 233
rect 23 226 27 231
rect 35 226 39 240
rect 85 244 87 246
rect 89 244 90 246
rect 23 222 39 226
rect 59 234 64 243
rect 50 233 64 234
rect 50 231 51 233
rect 53 231 54 233
rect 56 231 64 233
rect 50 230 64 231
rect 85 242 90 244
rect 159 250 171 251
rect 85 240 87 242
rect 89 240 90 242
rect 85 238 90 240
rect 58 225 71 226
rect 58 223 64 225
rect 66 223 71 225
rect 58 222 71 223
rect 23 219 27 222
rect -9 213 -7 215
rect -9 211 -5 213
rect -9 208 3 211
rect -9 206 -7 208
rect -5 206 3 208
rect -9 205 3 206
rect 15 213 27 219
rect 35 218 39 222
rect 35 216 40 218
rect 35 214 37 216
rect 39 214 40 216
rect 35 209 40 214
rect 67 216 71 222
rect 67 214 68 216
rect 70 214 71 216
rect 67 213 71 214
rect 85 215 89 238
rect 101 233 113 235
rect 101 231 104 233
rect 106 231 113 233
rect 101 229 113 231
rect 101 224 105 229
rect 101 222 102 224
rect 104 222 105 224
rect 101 221 105 222
rect 117 233 121 235
rect 119 231 121 233
rect 117 229 121 231
rect 142 234 147 243
rect 159 249 167 250
rect 159 247 160 249
rect 162 248 167 249
rect 169 248 171 250
rect 162 247 171 248
rect 159 245 171 247
rect 167 242 171 245
rect 169 240 171 242
rect 142 233 156 234
rect 142 231 144 233
rect 146 231 150 233
rect 152 231 156 233
rect 142 230 156 231
rect 117 227 118 229
rect 120 227 121 229
rect 117 219 121 227
rect 85 213 87 215
rect 35 207 37 209
rect 39 207 40 209
rect 35 205 40 207
rect 85 211 89 213
rect 85 208 97 211
rect 85 206 87 208
rect 89 206 97 208
rect 85 205 97 206
rect 109 213 121 219
rect 135 225 148 226
rect 135 223 140 225
rect 142 223 148 225
rect 135 222 148 223
rect 135 217 139 222
rect 167 218 171 240
rect 192 248 197 251
rect 192 246 193 248
rect 195 246 197 248
rect 211 249 229 250
rect 211 247 213 249
rect 215 247 229 249
rect 211 246 229 247
rect 192 242 197 246
rect 192 241 219 242
rect 192 239 194 241
rect 196 239 219 241
rect 192 238 219 239
rect 215 236 216 238
rect 218 236 219 238
rect 215 234 219 236
rect 192 233 209 234
rect 192 231 205 233
rect 207 231 209 233
rect 192 230 209 231
rect 192 228 197 230
rect 192 226 193 228
rect 195 226 197 228
rect 225 226 229 246
rect 192 221 197 226
rect 207 225 229 226
rect 207 223 226 225
rect 228 223 229 225
rect 207 221 208 223
rect 210 222 229 223
rect 210 221 213 222
rect 135 215 136 217
rect 138 215 139 217
rect 135 213 139 215
rect 166 216 171 218
rect 166 214 167 216
rect 169 214 171 216
rect 166 209 171 214
rect 207 216 213 221
rect 207 214 208 216
rect 210 214 213 216
rect 207 212 213 214
rect 166 207 167 209
rect 169 207 171 209
rect 166 205 171 207
rect -13 199 233 200
rect -25 197 4 199
rect 6 197 98 199
rect 100 197 233 199
rect -25 192 233 197
rect -25 163 -12 192
rect -25 158 238 163
rect -25 156 -2 158
rect 0 156 226 158
rect 228 156 238 158
rect -25 155 238 156
rect -25 9 -17 155
rect 88 148 93 150
rect 88 146 89 148
rect 91 146 93 148
rect 11 140 16 142
rect 11 138 13 140
rect 15 138 16 140
rect 3 126 7 134
rect 11 133 16 138
rect 35 133 39 134
rect 57 133 61 142
rect 88 141 93 146
rect 120 148 126 149
rect 120 146 122 148
rect 124 146 126 148
rect 88 139 89 141
rect 91 139 93 141
rect 88 137 93 139
rect 120 142 126 146
rect 135 148 140 150
rect 135 146 137 148
rect 139 146 140 148
rect 120 141 129 142
rect 120 139 122 141
rect 124 139 129 141
rect 120 138 129 139
rect 89 134 93 137
rect 11 131 13 133
rect 15 131 33 133
rect 35 132 70 133
rect 35 131 62 132
rect 11 130 62 131
rect 64 130 70 132
rect 11 129 70 130
rect -12 125 7 126
rect -12 123 -10 125
rect -8 124 24 125
rect -8 123 10 124
rect -12 122 10 123
rect 12 122 18 124
rect 20 122 24 124
rect -12 121 24 122
rect 35 117 39 129
rect 10 115 39 117
rect 10 113 13 115
rect 15 113 33 115
rect 35 113 39 115
rect 64 124 78 125
rect 64 122 72 124
rect 74 122 78 124
rect 64 121 78 122
rect 64 115 69 121
rect 89 132 113 134
rect 89 130 90 132
rect 92 130 113 132
rect 89 129 121 130
rect 10 108 16 113
rect 31 112 39 113
rect 64 113 66 115
rect 68 113 69 115
rect 64 112 69 113
rect 10 106 13 108
rect 15 106 16 108
rect 10 104 16 106
rect 89 115 93 129
rect 109 126 121 129
rect 117 124 121 126
rect 117 122 118 124
rect 120 122 121 124
rect 97 121 113 122
rect 97 119 98 121
rect 100 119 108 121
rect 110 119 113 121
rect 117 120 121 122
rect 97 118 113 119
rect 91 113 93 115
rect 89 110 93 113
rect 109 112 113 118
rect 81 107 93 110
rect 81 105 89 107
rect 91 105 93 107
rect 81 104 93 105
rect 125 110 129 138
rect 117 108 129 110
rect 112 107 129 108
rect 112 105 114 107
rect 116 105 129 107
rect 112 104 129 105
rect 135 141 140 146
rect 135 139 137 141
rect 139 139 140 141
rect 135 137 140 139
rect 135 126 139 137
rect 167 133 171 142
rect 187 133 191 134
rect 210 140 215 142
rect 210 138 211 140
rect 213 138 215 140
rect 210 133 215 138
rect 135 124 136 126
rect 138 124 139 126
rect 135 115 139 124
rect 158 132 191 133
rect 158 130 164 132
rect 166 131 191 132
rect 193 131 211 133
rect 213 131 215 133
rect 166 130 215 131
rect 158 129 215 130
rect 150 124 177 125
rect 150 122 154 124
rect 156 122 173 124
rect 175 122 177 124
rect 150 121 177 122
rect 135 113 137 115
rect 135 110 139 113
rect 135 107 147 110
rect 135 105 137 107
rect 139 105 147 107
rect 159 112 164 121
rect 187 117 191 129
rect 219 125 223 134
rect 202 124 227 125
rect 202 122 206 124
rect 208 122 214 124
rect 216 122 224 124
rect 226 122 227 124
rect 202 121 227 122
rect 187 115 216 117
rect 187 113 191 115
rect 193 113 211 115
rect 213 113 216 115
rect 187 112 195 113
rect 135 104 147 105
rect 210 108 216 113
rect 210 106 211 108
rect 213 106 216 108
rect 210 104 216 106
rect 246 99 255 256
rect -9 98 255 99
rect -9 96 42 98
rect 44 96 78 98
rect 80 96 104 98
rect 106 96 125 98
rect 127 96 148 98
rect 150 96 182 98
rect 184 96 253 98
rect -9 91 253 96
rect -9 73 3 91
rect -9 68 235 73
rect -9 66 42 68
rect 44 66 76 68
rect 78 66 99 68
rect 101 66 120 68
rect 122 66 146 68
rect 148 66 182 68
rect 184 66 235 68
rect -9 65 235 66
rect 10 58 16 60
rect 10 56 13 58
rect 15 56 16 58
rect 10 51 16 56
rect 79 59 91 60
rect 31 51 39 52
rect 10 49 13 51
rect 15 49 33 51
rect 35 49 39 51
rect 10 47 39 49
rect -1 42 24 43
rect -1 40 0 42
rect 2 40 10 42
rect 12 40 18 42
rect 20 40 24 42
rect -1 39 24 40
rect 3 30 7 39
rect 35 35 39 47
rect 62 43 67 52
rect 79 57 87 59
rect 89 57 91 59
rect 79 54 91 57
rect 87 51 91 54
rect 89 49 91 51
rect 49 42 76 43
rect 49 40 51 42
rect 53 40 70 42
rect 72 40 76 42
rect 49 39 76 40
rect 11 34 68 35
rect 11 33 60 34
rect 11 31 13 33
rect 15 31 33 33
rect 35 32 60 33
rect 62 32 68 34
rect 35 31 68 32
rect 87 40 91 49
rect 87 38 88 40
rect 90 38 91 40
rect 11 26 16 31
rect 11 24 13 26
rect 15 24 16 26
rect 11 22 16 24
rect 35 30 39 31
rect 55 22 59 31
rect 87 27 91 38
rect 86 25 91 27
rect 86 23 87 25
rect 89 23 91 25
rect 86 18 91 23
rect 97 59 114 60
rect 97 57 110 59
rect 112 57 114 59
rect 97 56 114 57
rect 97 54 109 56
rect 97 26 101 54
rect 133 59 145 60
rect 133 57 135 59
rect 137 57 145 59
rect 133 54 145 57
rect 113 46 117 52
rect 133 51 137 54
rect 133 49 135 51
rect 113 45 129 46
rect 105 42 109 44
rect 113 43 116 45
rect 118 43 126 45
rect 128 43 129 45
rect 113 42 129 43
rect 105 40 106 42
rect 108 40 109 42
rect 105 38 109 40
rect 105 35 117 38
rect 133 35 137 49
rect 210 58 216 60
rect 210 56 211 58
rect 213 56 216 58
rect 157 51 162 52
rect 157 49 158 51
rect 160 49 162 51
rect 187 51 195 52
rect 210 51 216 56
rect 105 34 134 35
rect 113 33 134 34
rect 136 33 137 35
rect 113 30 137 33
rect 157 43 162 49
rect 148 42 162 43
rect 148 40 152 42
rect 154 40 162 42
rect 148 39 162 40
rect 187 49 191 51
rect 193 49 211 51
rect 213 49 216 51
rect 187 47 216 49
rect 187 35 191 47
rect 202 42 238 43
rect 202 40 206 42
rect 208 40 214 42
rect 216 41 238 42
rect 216 40 234 41
rect 202 39 234 40
rect 236 39 238 41
rect 219 38 238 39
rect 156 34 215 35
rect 156 32 162 34
rect 164 33 215 34
rect 164 32 191 33
rect 156 31 191 32
rect 193 31 211 33
rect 213 31 215 33
rect 133 27 137 30
rect 97 25 106 26
rect 97 23 102 25
rect 104 23 106 25
rect 97 22 106 23
rect 86 16 87 18
rect 89 16 91 18
rect 86 14 91 16
rect 100 18 106 22
rect 133 25 138 27
rect 133 23 135 25
rect 137 23 138 25
rect 100 16 102 18
rect 104 16 106 18
rect 100 15 106 16
rect 133 18 138 23
rect 165 22 169 31
rect 187 30 191 31
rect 210 26 215 31
rect 219 30 223 38
rect 210 24 211 26
rect 213 24 215 26
rect 210 22 215 24
rect 133 16 135 18
rect 137 16 138 18
rect 133 14 138 16
rect -25 8 238 9
rect -25 6 -2 8
rect 0 6 226 8
rect 228 6 238 8
rect -25 1 238 6
<< alu2 >>
rect 85 268 239 274
rect 85 246 90 268
rect 85 244 87 246
rect 89 244 90 246
rect -9 238 -4 242
rect 85 238 90 244
rect 116 249 164 251
rect 116 247 160 249
rect 162 247 164 249
rect 116 245 164 247
rect 192 248 197 268
rect 192 246 193 248
rect 195 246 197 248
rect -9 236 -8 238
rect -6 236 -4 238
rect -9 234 -4 236
rect -9 232 -8 234
rect -6 232 -4 234
rect -9 228 -4 232
rect 50 233 58 234
rect 50 231 51 233
rect 53 231 58 233
rect 50 230 58 231
rect 7 227 11 228
rect 7 224 8 227
rect 10 224 11 227
rect 7 172 11 224
rect 54 186 58 230
rect 116 229 121 245
rect 192 244 197 246
rect 234 242 239 268
rect 234 237 264 242
rect 116 227 118 229
rect 120 227 121 229
rect 116 226 121 227
rect 143 233 148 234
rect 143 231 144 233
rect 146 231 148 233
rect 101 224 105 225
rect 101 222 102 224
rect 104 222 105 224
rect 101 221 105 222
rect 67 217 139 218
rect 67 216 136 217
rect 67 214 68 216
rect 70 215 136 216
rect 138 215 139 217
rect 70 214 139 215
rect 67 213 139 214
rect 54 184 55 186
rect 57 184 58 186
rect 54 183 58 184
rect 7 168 93 172
rect 89 132 93 168
rect 120 148 126 213
rect 143 178 148 231
rect 192 230 197 231
rect 192 226 193 230
rect 195 226 197 230
rect 192 225 197 226
rect 225 225 265 227
rect 225 223 226 225
rect 228 223 265 225
rect 225 222 265 223
rect 120 146 122 148
rect 124 146 126 148
rect 120 144 126 146
rect 135 172 148 178
rect 89 130 90 132
rect 92 130 93 132
rect 89 128 93 130
rect 135 127 140 172
rect 131 126 140 127
rect -12 125 -6 126
rect -12 123 -10 125
rect -8 123 -6 125
rect 131 124 136 126
rect 138 124 140 126
rect 131 123 140 124
rect 171 124 177 125
rect -12 91 -6 123
rect 171 122 173 124
rect 175 122 177 124
rect 96 121 101 122
rect 96 119 98 121
rect 100 119 101 121
rect 96 118 101 119
rect 64 115 69 116
rect 64 113 66 115
rect 68 113 69 115
rect 64 112 69 113
rect 126 111 138 112
rect 126 109 127 111
rect 129 109 138 111
rect 126 108 138 109
rect -12 86 55 91
rect -1 42 3 43
rect -1 40 0 42
rect 2 40 3 42
rect -1 39 3 40
rect 49 42 55 86
rect 125 45 130 46
rect 125 43 126 45
rect 128 43 130 45
rect 125 42 130 43
rect 49 40 51 42
rect 53 40 55 42
rect 49 39 55 40
rect 87 40 95 41
rect 87 38 88 40
rect 90 38 95 40
rect 87 37 95 38
rect 134 36 138 108
rect 171 78 177 122
rect 223 124 227 125
rect 223 122 224 124
rect 226 122 227 124
rect 223 121 227 122
rect 171 73 238 78
rect 157 51 162 52
rect 157 49 158 51
rect 160 49 162 51
rect 157 48 162 49
rect 232 41 238 73
rect 232 39 234 41
rect 236 39 238 41
rect 232 38 238 39
rect 133 35 138 36
rect 133 33 134 35
rect 136 33 138 35
rect 133 32 138 33
<< alu3 >>
rect -9 276 246 282
rect -9 238 -4 276
rect -9 236 -8 238
rect -6 236 -4 238
rect -9 228 -4 236
rect 173 231 179 276
rect 241 252 246 276
rect 241 248 264 252
rect 251 247 264 248
rect 173 230 197 231
rect 173 228 193 230
rect 195 228 197 230
rect 173 226 197 228
rect 101 224 105 225
rect 101 222 102 224
rect 104 222 105 224
rect 101 221 105 222
rect 54 186 130 187
rect 54 184 55 186
rect 57 184 130 186
rect 54 183 130 184
rect 96 121 101 122
rect 96 119 98 121
rect 100 119 101 121
rect 96 118 101 119
rect 64 115 69 116
rect 64 113 66 115
rect 68 113 69 115
rect 64 78 69 113
rect 126 112 130 183
rect 135 126 139 127
rect 135 124 136 126
rect 138 124 139 126
rect 135 123 139 124
rect 223 124 238 125
rect 223 122 224 124
rect 226 122 238 124
rect 223 121 238 122
rect 126 111 132 112
rect 126 109 127 111
rect 129 109 132 111
rect 126 108 132 109
rect 234 91 238 121
rect -12 73 69 78
rect 157 86 238 91
rect -12 43 -8 73
rect 157 51 162 86
rect 157 49 158 51
rect 160 49 162 51
rect 157 48 162 49
rect 125 45 130 46
rect 125 43 126 45
rect 128 43 130 45
rect -12 42 3 43
rect 125 42 130 43
rect -12 40 0 42
rect 2 40 3 42
rect -12 39 3 40
rect 87 40 95 41
rect 87 38 88 40
rect 90 38 95 40
rect 87 37 95 38
<< alu4 >>
rect 101 224 105 226
rect 101 222 102 224
rect 104 222 105 224
rect 101 181 105 222
rect 93 176 105 181
rect 93 122 97 176
rect 131 126 139 127
rect 131 124 136 126
rect 138 124 139 126
rect 131 123 139 124
rect 93 121 101 122
rect 93 119 98 121
rect 100 119 101 121
rect 93 118 101 119
rect 128 119 135 123
rect 93 111 99 118
rect 92 110 99 111
rect 92 45 98 110
rect 128 54 134 119
rect 127 53 134 54
rect 127 46 133 53
rect 91 41 98 45
rect 125 45 133 46
rect 125 43 126 45
rect 128 43 133 45
rect 125 42 133 43
rect 87 40 95 41
rect 87 38 88 40
rect 90 38 95 40
rect 87 37 95 38
<< ptie >>
rect 16 259 26 261
rect 16 257 20 259
rect 22 257 26 259
rect 110 259 120 261
rect 110 257 114 259
rect 116 257 120 259
rect 16 255 26 257
rect 110 255 120 257
rect 186 259 192 261
rect 186 257 188 259
rect 190 257 192 259
rect 186 246 192 257
rect 40 98 46 100
rect 40 96 42 98
rect 44 96 46 98
rect 40 94 46 96
rect 102 98 108 100
rect 102 96 104 98
rect 106 96 108 98
rect 102 94 108 96
rect 180 98 186 100
rect 180 96 182 98
rect 184 96 186 98
rect 180 94 186 96
rect 40 68 46 70
rect 40 66 42 68
rect 44 66 46 68
rect 40 64 46 66
rect 118 68 124 70
rect 118 66 120 68
rect 122 66 124 68
rect 118 64 124 66
rect 180 68 186 70
rect 180 66 182 68
rect 184 66 186 68
rect 180 64 186 66
<< ntie >>
rect -4 158 2 160
rect -4 156 -2 158
rect 0 156 2 158
rect 224 158 230 160
rect -4 154 2 156
rect 224 156 226 158
rect 228 156 230 158
rect 224 154 230 156
rect -4 8 2 10
rect -4 6 -2 8
rect 0 6 2 8
rect 224 8 230 10
rect -4 4 2 6
rect 224 6 226 8
rect 228 6 230 8
rect 224 4 230 6
<< nmos >>
rect -2 238 0 252
rect 8 243 10 251
rect 18 241 20 249
rect 42 238 44 252
rect 55 238 57 251
rect 62 238 64 251
rect 92 238 94 252
rect 102 243 104 251
rect 112 241 114 249
rect 142 238 144 251
rect 149 238 151 251
rect 162 238 164 252
rect 208 243 210 258
rect 218 243 220 258
rect 8 97 10 117
rect 18 97 20 117
rect 28 97 30 117
rect 38 108 40 117
rect 64 104 66 117
rect 71 104 73 117
rect 84 103 86 117
rect 108 106 110 114
rect 119 103 121 111
rect 142 103 144 117
rect 155 104 157 117
rect 162 104 164 117
rect 186 108 188 117
rect 196 97 198 117
rect 206 97 208 117
rect 216 97 218 117
rect 8 47 10 67
rect 18 47 20 67
rect 28 47 30 67
rect 38 47 40 56
rect 62 47 64 60
rect 69 47 71 60
rect 82 47 84 61
rect 105 53 107 61
rect 116 50 118 58
rect 140 47 142 61
rect 153 47 155 60
rect 160 47 162 60
rect 186 47 188 56
rect 196 47 198 67
rect 206 47 208 67
rect 216 47 218 67
<< pmos >>
rect -2 198 0 226
rect 11 198 13 226
rect 18 198 20 226
rect 42 198 44 226
rect 52 198 54 217
rect 62 198 64 217
rect 92 198 94 226
rect 105 198 107 226
rect 112 198 114 226
rect 142 198 144 217
rect 152 198 154 217
rect 162 198 164 226
rect 196 198 198 225
rect 203 198 205 225
rect 213 198 215 225
rect 220 198 222 225
rect 8 129 10 149
rect 18 129 20 157
rect 28 129 30 157
rect 38 129 40 157
rect 64 138 66 157
rect 74 138 76 157
rect 84 129 86 157
rect 110 129 112 157
rect 117 129 119 157
rect 142 129 144 157
rect 152 138 154 157
rect 162 138 164 157
rect 186 129 188 157
rect 196 129 198 157
rect 206 129 208 157
rect 216 129 218 149
rect 8 15 10 35
rect 18 7 20 35
rect 28 7 30 35
rect 38 7 40 35
rect 62 7 64 26
rect 72 7 74 26
rect 82 7 84 35
rect 107 7 109 35
rect 114 7 116 35
rect 140 7 142 35
rect 150 7 152 26
rect 160 7 162 26
rect 186 7 188 35
rect 196 7 198 35
rect 206 7 208 35
rect 216 15 218 35
<< polyct0 >>
rect 0 231 2 233
rect 44 231 46 233
rect 94 231 96 233
rect 160 231 162 233
rect 82 122 84 124
rect 144 122 146 124
rect 80 40 82 42
rect 142 40 144 42
<< polyct1 >>
rect 10 231 12 233
rect 23 231 25 233
rect 54 231 56 233
rect 194 239 196 241
rect 104 231 106 233
rect 117 231 119 233
rect 150 231 152 233
rect 64 223 66 225
rect 140 223 142 225
rect 216 236 218 238
rect 205 231 207 233
rect 62 130 64 132
rect 10 122 12 124
rect 18 122 20 124
rect 72 122 74 124
rect 164 130 166 132
rect 108 119 110 121
rect 118 122 120 124
rect 154 122 156 124
rect 206 122 208 124
rect 214 122 216 124
rect 10 40 12 42
rect 18 40 20 42
rect 70 40 72 42
rect 106 40 108 42
rect 116 43 118 45
rect 60 32 62 34
rect 152 40 154 42
rect 206 40 208 42
rect 214 40 216 42
rect 162 32 164 34
<< ndifct0 >>
rect 3 247 5 249
rect 13 245 15 247
rect 23 245 25 247
rect 67 247 69 249
rect 97 247 99 249
rect 107 245 109 247
rect 117 245 119 247
rect 137 247 139 249
rect 203 254 205 256
rect 203 247 205 249
rect 223 254 225 256
rect 2 106 4 108
rect 2 99 4 101
rect 23 106 25 108
rect 23 99 25 101
rect 43 110 45 112
rect 59 106 61 108
rect 103 108 105 110
rect 181 110 183 112
rect 167 106 169 108
rect 201 106 203 108
rect 201 99 203 101
rect 222 106 224 108
rect 222 99 224 101
rect 2 63 4 65
rect 2 56 4 58
rect 23 63 25 65
rect 23 56 25 58
rect 57 56 59 58
rect 43 52 45 54
rect 121 54 123 56
rect 165 56 167 58
rect 181 52 183 54
rect 201 63 203 65
rect 201 56 203 58
rect 222 63 224 65
rect 222 56 224 58
<< ndifct1 >>
rect 48 257 50 259
rect -7 247 -5 249
rect -7 240 -5 242
rect 37 248 39 250
rect 37 240 39 242
rect 87 247 89 249
rect 87 240 89 242
rect 156 257 158 259
rect 167 248 169 250
rect 213 247 215 249
rect 167 240 169 242
rect 13 113 15 115
rect 13 106 15 108
rect 33 113 35 115
rect 89 113 91 115
rect 89 105 91 107
rect 137 113 139 115
rect 114 105 116 107
rect 137 105 139 107
rect 191 113 193 115
rect 78 96 80 98
rect 125 96 127 98
rect 148 96 150 98
rect 211 113 213 115
rect 211 106 213 108
rect 13 56 15 58
rect 13 49 15 51
rect 76 66 78 68
rect 99 66 101 68
rect 146 66 148 68
rect 33 49 35 51
rect 87 57 89 59
rect 110 57 112 59
rect 87 49 89 51
rect 135 57 137 59
rect 135 49 137 51
rect 191 49 193 51
rect 211 56 213 58
rect 211 49 213 51
<< ntiect1 >>
rect -2 156 0 158
rect 226 156 228 158
rect -2 6 0 8
rect 226 6 228 8
<< ptiect1 >>
rect 20 257 22 259
rect 114 257 116 259
rect 188 257 190 259
rect 42 96 44 98
rect 104 96 106 98
rect 182 96 184 98
rect 42 66 44 68
rect 120 66 122 68
rect 182 66 184 68
<< pdifct0 >>
rect 23 206 25 208
rect 47 207 49 209
rect 47 200 49 202
rect 57 213 59 215
rect 57 206 59 208
rect 67 207 69 209
rect 67 200 69 202
rect 117 206 119 208
rect 137 207 139 209
rect 137 200 139 202
rect 147 213 149 215
rect 147 206 149 208
rect 157 207 159 209
rect 157 200 159 202
rect 191 207 193 209
rect 191 200 193 202
rect 225 207 227 209
rect 225 200 227 202
rect 3 145 5 147
rect 3 138 5 140
rect 23 153 25 155
rect 23 145 25 147
rect 33 138 35 140
rect 43 153 45 155
rect 43 146 45 148
rect 59 153 61 155
rect 59 146 61 148
rect 69 147 71 149
rect 69 140 71 142
rect 79 153 81 155
rect 79 146 81 148
rect 103 153 105 155
rect 103 146 105 148
rect 147 153 149 155
rect 147 146 149 148
rect 157 147 159 149
rect 157 140 159 142
rect 167 153 169 155
rect 167 146 169 148
rect 181 153 183 155
rect 181 146 183 148
rect 191 138 193 140
rect 201 153 203 155
rect 201 145 203 147
rect 221 145 223 147
rect 221 138 223 140
rect 3 24 5 26
rect 3 17 5 19
rect 23 17 25 19
rect 23 9 25 11
rect 33 24 35 26
rect 43 16 45 18
rect 43 9 45 11
rect 57 16 59 18
rect 57 9 59 11
rect 67 22 69 24
rect 67 15 69 17
rect 77 16 79 18
rect 77 9 79 11
rect 121 16 123 18
rect 121 9 123 11
rect 145 16 147 18
rect 145 9 147 11
rect 155 22 157 24
rect 155 15 157 17
rect 165 16 167 18
rect 165 9 167 11
rect 181 16 183 18
rect 181 9 183 11
rect 191 24 193 26
rect 201 17 203 19
rect 201 9 203 11
rect 221 24 223 26
rect 221 17 223 19
<< pdifct1 >>
rect -7 213 -5 215
rect -7 206 -5 208
rect 4 197 6 199
rect 37 214 39 216
rect 37 207 39 209
rect 87 213 89 215
rect 87 206 89 208
rect 98 197 100 199
rect 167 214 169 216
rect 167 207 169 209
rect 208 221 210 223
rect 208 214 210 216
rect 13 138 15 140
rect 13 131 15 133
rect 33 131 35 133
rect 89 146 91 148
rect 89 139 91 141
rect 122 146 124 148
rect 122 139 124 141
rect 137 146 139 148
rect 137 139 139 141
rect 191 131 193 133
rect 211 138 213 140
rect 211 131 213 133
rect 13 31 15 33
rect 13 24 15 26
rect 33 31 35 33
rect 87 23 89 25
rect 87 16 89 18
rect 102 23 104 25
rect 102 16 104 18
rect 135 23 137 25
rect 135 16 137 18
rect 191 31 193 33
rect 211 31 213 33
rect 211 24 213 26
<< alu0 >>
rect 1 249 7 256
rect 1 247 3 249
rect 5 247 7 249
rect 1 246 7 247
rect 12 247 16 249
rect 12 245 13 247
rect 15 245 16 247
rect 12 243 16 245
rect 21 247 27 256
rect 21 245 23 247
rect 25 245 27 247
rect 21 244 27 245
rect 51 249 71 250
rect 51 247 67 249
rect 69 247 71 249
rect 51 246 71 247
rect 95 249 101 256
rect 95 247 97 249
rect 99 247 101 249
rect 95 246 101 247
rect 106 247 110 249
rect -1 239 16 243
rect -1 233 3 239
rect -1 231 0 233
rect 2 231 3 233
rect -1 218 3 231
rect 22 219 23 235
rect 39 238 40 245
rect 51 242 55 246
rect 43 238 55 242
rect 43 233 47 238
rect 43 231 44 233
rect 46 231 47 233
rect 43 226 47 231
rect 106 245 107 247
rect 109 245 110 247
rect 106 243 110 245
rect 115 247 121 256
rect 201 254 203 256
rect 205 254 207 256
rect 115 245 117 247
rect 119 245 121 247
rect 135 249 155 250
rect 135 247 137 249
rect 139 247 155 249
rect 135 246 155 247
rect 115 244 121 245
rect 93 239 110 243
rect 43 222 51 226
rect -5 211 -4 217
rect -1 214 11 218
rect 7 209 11 214
rect 47 218 51 222
rect 47 215 61 218
rect 47 214 57 215
rect 55 213 57 214
rect 59 213 61 215
rect 93 233 97 239
rect 93 231 94 233
rect 96 231 97 233
rect 93 218 97 231
rect 116 219 117 235
rect 151 242 155 246
rect 151 238 163 242
rect 166 238 167 245
rect 159 233 163 238
rect 159 231 160 233
rect 162 231 163 233
rect 159 226 163 231
rect 7 208 27 209
rect 7 206 23 208
rect 25 206 27 208
rect 7 205 27 206
rect 45 209 51 210
rect 45 207 47 209
rect 49 207 51 209
rect 45 202 51 207
rect 55 208 61 213
rect 89 211 90 217
rect 93 214 105 218
rect 55 206 57 208
rect 59 206 61 208
rect 55 205 61 206
rect 65 209 71 210
rect 65 207 67 209
rect 69 207 71 209
rect 45 200 47 202
rect 49 200 51 202
rect 65 202 71 207
rect 101 209 105 214
rect 155 222 163 226
rect 155 218 159 222
rect 201 249 207 254
rect 221 254 223 256
rect 225 254 227 256
rect 221 253 227 254
rect 201 247 203 249
rect 205 247 207 249
rect 201 246 207 247
rect 145 215 159 218
rect 145 213 147 215
rect 149 214 159 215
rect 149 213 151 214
rect 135 209 141 210
rect 101 208 121 209
rect 101 206 117 208
rect 119 206 121 208
rect 101 205 121 206
rect 135 207 137 209
rect 139 207 141 209
rect 65 200 67 202
rect 69 200 71 202
rect 135 202 141 207
rect 145 208 151 213
rect 145 206 147 208
rect 149 206 151 208
rect 145 205 151 206
rect 155 209 161 210
rect 155 207 157 209
rect 159 207 161 209
rect 135 200 137 202
rect 139 200 141 202
rect 155 202 161 207
rect 189 209 195 210
rect 189 207 191 209
rect 193 207 195 209
rect 155 200 157 202
rect 159 200 161 202
rect 189 202 195 207
rect 189 200 191 202
rect 193 200 195 202
rect 223 209 229 210
rect 223 207 225 209
rect 227 207 229 209
rect 223 202 229 207
rect 223 200 225 202
rect 227 200 229 202
rect 1 147 7 155
rect 1 145 3 147
rect 5 145 7 147
rect 1 140 7 145
rect 22 153 23 155
rect 25 153 26 155
rect 22 147 26 153
rect 22 145 23 147
rect 25 145 26 147
rect 41 153 43 155
rect 45 153 47 155
rect 41 148 47 153
rect 41 146 43 148
rect 45 146 47 148
rect 41 145 47 146
rect 57 153 59 155
rect 61 153 63 155
rect 57 148 63 153
rect 77 153 79 155
rect 81 153 83 155
rect 57 146 59 148
rect 61 146 63 148
rect 57 145 63 146
rect 67 149 73 150
rect 67 147 69 149
rect 71 147 73 149
rect 22 143 26 145
rect 67 142 73 147
rect 77 148 83 153
rect 102 153 103 155
rect 105 153 106 155
rect 77 146 79 148
rect 81 146 83 148
rect 77 145 83 146
rect 1 138 3 140
rect 5 138 7 140
rect 1 137 7 138
rect 32 140 36 142
rect 32 138 33 140
rect 35 138 36 140
rect 32 134 36 138
rect 32 133 35 134
rect 67 140 69 142
rect 71 141 73 142
rect 102 148 106 153
rect 145 153 147 155
rect 149 153 151 155
rect 102 146 103 148
rect 105 146 106 148
rect 102 144 106 146
rect 71 140 81 141
rect 67 137 81 140
rect 77 133 81 137
rect 77 129 85 133
rect 81 124 85 129
rect 81 122 82 124
rect 84 122 85 124
rect 81 117 85 122
rect 0 108 6 109
rect 0 106 2 108
rect 4 106 6 108
rect 0 101 6 106
rect 42 112 46 114
rect 73 113 85 117
rect 42 110 43 112
rect 45 110 46 112
rect 21 108 27 109
rect 21 106 23 108
rect 25 106 27 108
rect 0 99 2 101
rect 4 99 6 101
rect 21 101 27 106
rect 21 99 23 101
rect 25 99 27 101
rect 42 99 46 110
rect 73 109 77 113
rect 88 110 89 117
rect 57 108 77 109
rect 57 106 59 108
rect 61 106 77 108
rect 57 105 77 106
rect 102 110 106 112
rect 102 108 103 110
rect 105 108 106 110
rect 102 99 106 108
rect 145 148 151 153
rect 165 153 167 155
rect 169 153 171 155
rect 145 146 147 148
rect 149 146 151 148
rect 145 145 151 146
rect 155 149 161 150
rect 155 147 157 149
rect 159 147 161 149
rect 155 142 161 147
rect 165 148 171 153
rect 165 146 167 148
rect 169 146 171 148
rect 165 145 171 146
rect 179 153 181 155
rect 183 153 185 155
rect 179 148 185 153
rect 179 146 181 148
rect 183 146 185 148
rect 179 145 185 146
rect 200 153 201 155
rect 203 153 204 155
rect 200 147 204 153
rect 200 145 201 147
rect 203 145 204 147
rect 200 143 204 145
rect 219 147 225 155
rect 219 145 221 147
rect 223 145 225 147
rect 155 141 157 142
rect 147 140 157 141
rect 159 140 161 142
rect 147 137 161 140
rect 147 133 151 137
rect 190 140 194 142
rect 190 138 191 140
rect 193 138 194 140
rect 190 134 194 138
rect 191 133 194 134
rect 219 140 225 145
rect 219 138 221 140
rect 223 138 225 140
rect 219 137 225 138
rect 143 129 151 133
rect 143 124 147 129
rect 143 122 144 124
rect 146 122 147 124
rect 143 117 147 122
rect 139 110 140 117
rect 143 113 155 117
rect 151 109 155 113
rect 180 112 184 114
rect 180 110 181 112
rect 183 110 184 112
rect 151 108 171 109
rect 151 106 167 108
rect 169 106 171 108
rect 151 105 171 106
rect 180 99 184 110
rect 199 108 205 109
rect 199 106 201 108
rect 203 106 205 108
rect 199 101 205 106
rect 220 108 226 109
rect 220 106 222 108
rect 224 106 226 108
rect 199 99 201 101
rect 203 99 205 101
rect 220 101 226 106
rect 220 99 222 101
rect 224 99 226 101
rect 0 63 2 65
rect 4 63 6 65
rect 0 58 6 63
rect 21 63 23 65
rect 25 63 27 65
rect 0 56 2 58
rect 4 56 6 58
rect 0 55 6 56
rect 21 58 27 63
rect 21 56 23 58
rect 25 56 27 58
rect 21 55 27 56
rect 42 54 46 65
rect 55 58 75 59
rect 55 56 57 58
rect 59 56 75 58
rect 55 55 75 56
rect 42 52 43 54
rect 45 52 46 54
rect 42 50 46 52
rect 71 51 75 55
rect 71 47 83 51
rect 86 47 87 54
rect 79 42 83 47
rect 79 40 80 42
rect 82 40 83 42
rect 79 35 83 40
rect 75 31 83 35
rect 1 26 7 27
rect 1 24 3 26
rect 5 24 7 26
rect 1 19 7 24
rect 32 30 35 31
rect 32 26 36 30
rect 32 24 33 26
rect 35 24 36 26
rect 32 22 36 24
rect 75 27 79 31
rect 65 24 79 27
rect 65 22 67 24
rect 69 23 79 24
rect 69 22 71 23
rect 1 17 3 19
rect 5 17 7 19
rect 1 9 7 17
rect 22 19 26 21
rect 22 17 23 19
rect 25 17 26 19
rect 22 11 26 17
rect 22 9 23 11
rect 25 9 26 11
rect 41 18 47 19
rect 41 16 43 18
rect 45 16 47 18
rect 41 11 47 16
rect 41 9 43 11
rect 45 9 47 11
rect 55 18 61 19
rect 55 16 57 18
rect 59 16 61 18
rect 55 11 61 16
rect 65 17 71 22
rect 65 15 67 17
rect 69 15 71 17
rect 65 14 71 15
rect 75 18 81 19
rect 75 16 77 18
rect 79 16 81 18
rect 55 9 57 11
rect 59 9 61 11
rect 75 11 81 16
rect 120 56 124 65
rect 120 54 121 56
rect 123 54 124 56
rect 120 52 124 54
rect 149 58 169 59
rect 149 56 165 58
rect 167 56 169 58
rect 149 55 169 56
rect 137 47 138 54
rect 149 51 153 55
rect 180 54 184 65
rect 199 63 201 65
rect 203 63 205 65
rect 199 58 205 63
rect 220 63 222 65
rect 224 63 226 65
rect 199 56 201 58
rect 203 56 205 58
rect 199 55 205 56
rect 180 52 181 54
rect 183 52 184 54
rect 141 47 153 51
rect 180 50 184 52
rect 220 58 226 63
rect 220 56 222 58
rect 224 56 226 58
rect 220 55 226 56
rect 141 42 145 47
rect 141 40 142 42
rect 144 40 145 42
rect 141 35 145 40
rect 141 31 149 35
rect 145 27 149 31
rect 145 24 159 27
rect 145 23 155 24
rect 120 18 124 20
rect 120 16 121 18
rect 123 16 124 18
rect 75 9 77 11
rect 79 9 81 11
rect 120 11 124 16
rect 153 22 155 23
rect 157 22 159 24
rect 191 30 194 31
rect 190 26 194 30
rect 190 24 191 26
rect 193 24 194 26
rect 190 22 194 24
rect 219 26 225 27
rect 219 24 221 26
rect 223 24 225 26
rect 143 18 149 19
rect 143 16 145 18
rect 147 16 149 18
rect 120 9 121 11
rect 123 9 124 11
rect 143 11 149 16
rect 153 17 159 22
rect 200 19 204 21
rect 153 15 155 17
rect 157 15 159 17
rect 153 14 159 15
rect 163 18 169 19
rect 163 16 165 18
rect 167 16 169 18
rect 143 9 145 11
rect 147 9 149 11
rect 163 11 169 16
rect 163 9 165 11
rect 167 9 169 11
rect 179 18 185 19
rect 179 16 181 18
rect 183 16 185 18
rect 179 11 185 16
rect 179 9 181 11
rect 183 9 185 11
rect 200 17 201 19
rect 203 17 204 19
rect 200 11 204 17
rect 200 9 201 11
rect 203 9 204 11
rect 219 19 225 24
rect 219 17 221 19
rect 223 17 225 19
rect 219 9 225 17
<< via1 >>
rect -8 232 -6 234
rect 8 224 10 227
rect 87 244 89 246
rect 51 231 53 233
rect 68 214 70 216
rect 102 222 104 224
rect 160 247 162 249
rect 144 231 146 233
rect 118 227 120 229
rect 193 246 195 248
rect 193 226 195 228
rect 226 223 228 225
rect 136 215 138 217
rect 122 146 124 148
rect -10 123 -8 125
rect 90 130 92 132
rect 66 113 68 115
rect 98 119 100 121
rect 136 124 138 126
rect 173 122 175 124
rect 224 122 226 124
rect 0 40 2 42
rect 51 40 53 42
rect 88 38 90 40
rect 126 43 128 45
rect 158 49 160 51
rect 134 33 136 35
rect 234 39 236 41
<< via2 >>
rect -8 236 -6 238
rect 102 222 104 224
rect 55 184 57 186
rect 193 228 195 230
rect 136 124 138 126
rect 98 119 100 121
rect 66 113 68 115
rect 127 109 129 111
rect 0 40 2 42
rect 126 43 128 45
rect 88 38 90 40
rect 224 122 226 124
rect 158 49 160 51
<< via3 >>
rect 102 222 104 224
rect 98 119 100 121
rect 136 124 138 126
rect 126 43 128 45
rect 88 38 90 40
<< labels >>
rlabel alu1 39 94 39 95 1 vss
rlabel alu1 2 122 2 122 1 A0
rlabel alu1 37 119 37 119 1 neg_A0
rlabel alu1 67 119 67 119 1 B0
rlabel alu1 5 40 5 40 1 B0
rlabel alu1 37 43 37 43 1 neg_B0
rlabel alu1 126 119 126 119 7 Equal_a0_b0
rlabel alu1 95 131 95 131 1 Lt_a0_b0
rlabel alu4 94 44 94 44 1 Gt_a0_b0
rlabel alu1 133 36 137 40 5 Lt_A1_B1
rlabel alu1 99 43 99 43 3 Equal_A1_B1
rlabel alu1 137 122 137 122 5 Gt_A1_B1
rlabel alu1 190 121 190 121 5 neg_B1
rlabel alu1 221 122 221 122 5 B1
rlabel alu1 189 43 189 43 5 neg_A1
rlabel alu1 222 41 222 41 5 A1
rlabel alu1 187 69 187 70 5 vss
rlabel nwell 95 1 234 9 5 vdd
rlabel nwell -8 155 131 163 1 vdd
rlabel alu1 153 260 153 260 2 vss
rlabel alu1 153 196 153 196 2 vdd
rlabel alu1 169 229 169 229 1 GT_a_B_cas1
rlabel alu1 103 260 103 260 8 vss
rlabel alu1 103 196 103 196 8 vdd
rlabel alu1 86 228 86 228 1 2bit_greater
rlabel alu1 53 260 53 260 8 vss
rlabel alu1 53 196 53 196 8 vdd
rlabel alu1 9 260 9 260 8 vss
rlabel alu1 9 196 9 196 8 vdd
rlabel alu1 -8 227 -8 227 1 2bit_less
rlabel alu1 34 224 34 224 1 2bit_less_case1
rlabel alu1 207 260 207 260 2 vss
rlabel alu1 207 196 207 196 2 vdd
rlabel alu1 227 235 227 235 1 2bit_equal
rlabel alu2 248 239 248 239 7 2bit_greater
rlabel alu3 247 250 247 250 7 2bit_less
rlabel alu2 248 224 248 224 7 2bit_equal
<< end >>
